module cs_data(

output [229:0] w0,
output [229:0] w1,
output [229:0] w2,
output [229:0] w3,
output [229:0] w4,
output [229:0] w5,
output [229:0] w6,
output [229:0] w7,
output [229:0] w8,
output [229:0] w9,
output [229:0] w10,
output [229:0] w11,
output [229:0] w12,
output [229:0] w13,
output [229:0] w14,
output [229:0] w15,
output [229:0] w16,
output [229:0] w17,
output [229:0] w18,
output [229:0] w19,
output [229:0] w20,
output [229:0] w21,
output [229:0] w22,
output [229:0] w23,
output [229:0] w24,
output [229:0] w25,
output [229:0] w26,
output [229:0] w27,
output [229:0] w28,
output [229:0] w29,
output [229:0] w30,
output [229:0] w31,
output [229:0] w32,
output [229:0] w33,
output [229:0] w34,
output [229:0] w35,
output [229:0] w36,
output [229:0] w37,
output [229:0] w38,
output [229:0] w39,
output [229:0] w40,
output [229:0] w41,
output [229:0] w42,
output [229:0] w43,
output [229:0] w44,
output [229:0] w45,
output [229:0] w46,
output [229:0] w47,
output [229:0] w48,
output [229:0] w49,
output [229:0] w50,
output [229:0] w51,
output [229:0] w52,
output [229:0] w53,
output [229:0] w54,
output [229:0] w55,
output [229:0] w56,
output [229:0] w57,
output [229:0] w58,
output [229:0] w59,
output [229:0] w60,
output [229:0] w61,
output [229:0] w62,
output [229:0] w63,
output [229:0] w64,
output [229:0] w65,
output [229:0] w66,
output [229:0] w67,
output [229:0] w68,
output [229:0] w69,
output [229:0] w70,
output [229:0] w71,
output [229:0] w72,
output [229:0] w73,
output [229:0] w74,
output [229:0] w75,
output [229:0] w76,
output [229:0] w77,
output [229:0] w78,
output [229:0] w79,
output [229:0] w80,
output [229:0] w81,
output [229:0] w82,
output [229:0] w83,
output [229:0] w84,
output [229:0] w85,
output [229:0] w86,
output [229:0] w87,
output [229:0] w88,
output [229:0] w89,
output [229:0] w90,
output [229:0] w91,
output [229:0] w92,
output [229:0] w93,
output [229:0] w94,
output [229:0] w95,
output [229:0] w96,
output [229:0] w97,
output [229:0] w98,
output [229:0] w99,
output [229:0] w100,
output [229:0] w101,
output [229:0] w102,
output [229:0] w103,
output [229:0] w104,
output [229:0] w105,
output [229:0] w106,
output [229:0] w107,
output [229:0] w108,
output [229:0] w109,
output [229:0] w110,
output [229:0] w111,
output [229:0] w112,
output [229:0] w113,
output [229:0] w114,
output [229:0] w115,
output [229:0] w116,
output [229:0] w117,
output [229:0] w118,
output [229:0] w119,
output [229:0] w120,
output [229:0] w121,
output [229:0] w122,
output [229:0] w123,
output [229:0] w124,
output [229:0] w125,
output [229:0] w126,
output [229:0] w127,
output [229:0] w128,
output [229:0] w129,
output [229:0] w130,
output [229:0] w131,
output [229:0] w132,
output [229:0] w133,
output [229:0] w134,
output [229:0] w135,
output [229:0] w136,
output [229:0] w137,
output [229:0] w138,
output [229:0] w139);
assign w0 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_1_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w1 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_1_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w2 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_1_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w3 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_1_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w4 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_1_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w5 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_1_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w6 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_1_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w7 = {1'b1, 1'b1, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_1_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w8 = {1'b1, 1'b1, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_1_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w9 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00000, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0010, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w10 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00000, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0010, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w11 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00000, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0010, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w12 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00000, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0010, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w13 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00000, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0010, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w14 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00000, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0010, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w15 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00000, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0010, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w16 = {1'b1, 1'b1, 1'b0, 8'h00, 5'b00000, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0010, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w17 = {1'b1, 1'b1, 1'b0, 8'h00, 5'b00000, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0010, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w18 = {1'b1, 1'b1, 1'b1, 8'hBC, 5'b00010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_0100, 18'b000000000_0_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w19 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0000_1000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b1, 1'b0, 1'b1, 2'b10, 2'b10, 3'b000, 3'b100, 3'b101, 3'b000, 3'b010, 3'b000, 3'b000, 3'b000, 13'h0400, 13'h1000, 13'h0400, 13'h0002, 13'h0400, 13'h0001, 13'h0100, 13'h0002, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 2'b01, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w20 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0100_0000_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b1, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0400, 13'h0008, 13'h0400, 13'h0001, 13'h0200, 13'h0008, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 2'b10, 2'b01, 2'b01, 1'b0, 4'b0000};
assign w21 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_1000_0000_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b1, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b100, 3'b101, 3'b000, 3'b010, 3'b000, 3'b000, 3'b000, 13'h1000, 13'h1000, 13'h0800, 13'h0010, 13'h0001, 13'h0001, 13'h0100, 13'h0010, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 2'b01, 2'b00, 2'b00, 1'b0, 4'b1000};
assign w22 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00101, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0001_0000, 18'b000000000_0_1_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w23 = {1'b1, 1'b1, 1'b1, 8'h42, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0100_0000, 18'b000000000__0_00_0_0_0_0_0, 2'b01, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w24 = {1'b1, 1'b0, 1'b1, 8'hB0, 5'b00111, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_1000_0000, 18'b000000000_1_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0008, 13'h0001, 13'h0100, 13'h0001, 13'h0008, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w25 = {1'b1, 1'b0, 1'b1, 8'hB1, 5'b00111, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_1000_0000, 18'b000000000_1_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0008, 13'h0001, 13'h0100, 13'h0001, 13'h0008, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w26 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b01000, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0001_0000_0000, 18'b000000000_0_0_00_1_1_1_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w27 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0010_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w28 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0100_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w29 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_1000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b11, 1'b0, 1'b1, 1'b0, 1'b1, 2'b00, 2'b00, 3'b000, 3'b100, 3'b101, 3'b000, 3'b010, 3'b000, 3'b000, 3'b000, 13'h0400, 13'h1000, 13'h0001, 13'h0001, 13'h0400, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w30 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_1000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b10, 1'b0, 1'b1, 1'b0, 1'b1, 2'b00, 2'b00, 3'b000, 3'b100, 3'b101, 3'b000, 3'b010, 3'b000, 3'b000, 3'b000, 13'h0400, 13'h1000, 13'h0001, 13'h0001, 13'h0400, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w31 = {1'b0, 1'b0, 1'b1, 8'h87, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_1000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b11, 1'b0, 1'b1, 1'b0, 1'b1, 2'b10, 2'b10, 3'b000, 3'b100, 3'b101, 3'b000, 3'b010, 3'b000, 3'b000, 3'b000, 13'h0400, 13'h1000, 13'h0001, 13'h0001, 13'h0400, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w32 = {1'b0, 1'b0, 1'b1, 8'h85, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_1000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b10, 1'b0, 1'b1, 1'b0, 1'b1, 2'b10, 2'b10, 3'b000, 3'b100, 3'b101, 3'b000, 3'b010, 3'b000, 3'b000, 3'b000, 13'h0400, 13'h1000, 13'h0001, 13'h0001, 13'h0400, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w33 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_1000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b1, 1'b0, 1'b1, 2'b00, 2'b00, 3'b000, 3'b100, 3'b101, 3'b000, 3'b010, 3'b000, 3'b000, 3'b000, 13'h0400, 13'h1000, 13'h0001, 13'h0001, 13'h0400, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w34 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_1000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b1, 1'b0, 1'b1, 2'b10, 2'b10, 3'b000, 3'b100, 3'b101, 3'b000, 3'b010, 3'b000, 3'b000, 3'b000, 13'h0400, 13'h1000, 13'h0001, 13'h0001, 13'h0400, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w35 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0100_0000_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b1, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0400, 13'h0008, 13'h0400, 13'h0001, 13'h0200, 13'h0008, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 2'b10, 2'b01, 2'b01, 1'b0, 4'b0000};
assign w36 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0001_0000_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b1, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b100, 3'b101, 3'b000, 3'b010, 3'b000, 3'b000, 3'b000, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 2'b10, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w37 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w38 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w39 = {1'b1, 1'b1, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w40 = {1'b1, 1'b1, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w41 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b01, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0040, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b1, 4'b0000};
assign w42 = {1'b1, 1'b1, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b01, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0040, 13'h0100, 13'h0001, 13'h0001, 13'h0040, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b1, 4'b0000};
assign w43 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'd0, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w44 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'd1, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w45 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'd2, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w46 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'd3, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w47 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'd4, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w48 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'd5, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w49 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'd6, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w50 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'd7, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w51 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'd0, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w52 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'd1, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w53 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'd2, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w54 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'd3, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w55 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'd4, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w56 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'd5, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w57 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'd6, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w58 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'd7, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w59 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w60 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0010_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w61 = {1'b1, 1'b1, 1'b1, 8'h6F, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0100_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b11, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w62 = {1'b1, 1'b0, 1'b1, 8'h7F, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0100_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b11, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w63 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_1000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b110, 3'b001, 3'b111, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0002, 13'h0008, 13'h0004, 13'h0200, 13'h0002, 13'h0008, 13'h0004, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 2'b10, 2'b01, 2'b00, 1'b0, 4'b0001};
assign w64 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_1000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b110, 3'b001, 3'b111, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0002, 13'h0008, 13'h0004, 13'h0200, 13'h0002, 13'h0008, 13'h0004, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 2'b10, 2'b01, 2'b00, 1'b0, 4'b0100};
assign w65 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b01001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0001_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w66 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b01001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0001_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w67 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b01010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0010_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w68 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b01010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0010_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 13'h0001, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w69 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b01010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0010_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w70 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b01010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0010_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w71 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b01010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0010_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 13'h0100, 13'h1000, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w72 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b01010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0010_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w73 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b01010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0010_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w74 = {1'b1, 1'b1, 1'b0, 8'h00, 5'b01010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0010_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w75 = {1'b1, 1'b1, 1'b0, 8'h00, 5'b01010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0010_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w76 = {1'b1, 1'b1, 1'b1, 8'hFD, 5'b01011, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0100_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b11, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w77 = {1'b1, 1'b1, 1'b1, 8'hFE, 5'b01100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_1000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b11, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w78 = {1'b1, 1'b1, 1'b1, 8'h63, 5'b01101, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0001_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b11, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w79 = {1'b1, 1'b1, 1'b1, 8'h6B, 5'b01110, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0010_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b11, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w80 = {1'b1, 1'b1, 1'b1, 8'h68, 5'b01111, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0100_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b11, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w81 = {1'b1, 1'b1, 1'b1, 8'h69, 5'b10000, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_1000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b11, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b00, 2'b10, 1'b0, 4'b0000};
assign w82 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0100, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b01, 2'b10, 2'b01, 1'b0, 4'b0000};
assign w83 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd0, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w84 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd1, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w85 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd2, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w86 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd3, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w87 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd4, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w88 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd5, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w89 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd6, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w90 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd7, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w91 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b011, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0010, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w92 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b000, 3'b010, 3'b000, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0010, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w93 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0010, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w94 = {1'b0, 1'b0, 1'b1, 8'hA1, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0010, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w95 = {1'b0, 1'b0, 1'b1, 8'hA9, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0001_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b101, 3'b010, 3'b101, 3'b000, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 13'h0010, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w96 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b10, 2'b01, 2'b01, 1'b0, 4'b0000};
assign w97 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd0, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w98 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd1, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w99 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd2, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w100 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd3, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w101 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd4, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w102 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd5, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w103 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd6, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w104 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd7, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w105 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h1000, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w106 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b10, 2'b10, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b101, 3'b000, 13'h1000, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w107 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b000, 3'b010, 3'b101, 3'b000, 13'h0010, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w108 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 13'h0010, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w109 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 3'b011, 3'b000, 13'h0010, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w110 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b000, 3'b010, 3'b000, 3'b000, 13'h0010, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w111 = {1'b0, 1'b0, 1'b1, 8'hA0, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b100, 3'b010, 3'b100, 3'b000, 13'h0010, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w112 = {1'b0, 1'b0, 1'b1, 8'hA8, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0100_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b101, 3'b010, 3'b101, 3'b000, 13'h0010, 13'h0001, 13'h0001, 13'h0008, 13'h0200, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 2'b00, 2'b01, 2'b00, 1'b0, 4'b0000};
assign w113 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0001_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b1, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 13'h0001, 3'b000, 13'h0200, 13'h1000, 13'h0001, 13'h0008, 13'h0400, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w114 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b1_0000_0000_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b1, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 13'h0001, 3'b000, 13'h0200, 13'h1000, 13'h0001, 13'h0008, 13'h0800, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b1000};
assign w115 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b0_0000_0001_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b1, 1'b0, 1'b1, 2'b01, 2'b00, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 13'h0001, 3'b000, 13'h0200, 13'h1000, 13'h0001, 13'h0008, 13'h0400, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b0000};
assign w116 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00100, 3'b000, 1'b0, 1'b0, 37'b1_0000_0000_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b1, 1'b0, 1'b1, 2'b01, 2'b10, 3'b000, 3'b000, 3'b101, 3'b100, 3'b011, 3'b010, 13'h0001, 3'b000, 13'h0200, 13'h1000, 13'h0001, 13'h0008, 13'h0800, 13'h0001, 13'h0001, 13'h0008, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 2'b00, 1'b0, 4'b1000};
assign w117 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b10010, 3'b000, 1'b0, 1'b1, 37'b0_0000_0010_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b001, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w118 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b10010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0010_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b001, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w119 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b10010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0010_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'b001, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w120 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b10010, 3'b000, 1'b0, 1'b1, 37'b0_0000_0010_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b001, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w121 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b10010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0010_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b001, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w122 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b10010, 3'b000, 1'b0, 1'b0, 37'b0_0000_0010_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b10, 3'b001, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w123 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b10001, 3'b000, 1'b0, 1'b1, 37'b0_0000_0100_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b001, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w124 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b10001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0100_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b001, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w125 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b10001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0100_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b00, 3'b001, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w126 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b10001, 3'b000, 1'b0, 1'b1, 37'b0_0000_0100_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b001, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w127 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b10001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0100_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b001, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w128 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b10001, 3'b000, 1'b0, 1'b0, 37'b0_0000_0100_0000_0000_0000_0000_0000_0000_0000, 18'b000000000_1_0_00_1_1_0_1_1, 2'b00, 1'b0, 1'b0, 1'b0, 1'b1, 2'b00, 2'b10, 3'b001, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w129 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00110, 3'b000, 1'b0, 1'b0, 37'b0_0000_0000_0000_0000_0000_0000_0000_0010_0000, 18'b000000000_0_1_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 13'h0001, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w130 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0010_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd0, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w131 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0010_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd1, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w132 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0010_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd2, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w133 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0010_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd3, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w134 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0010_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd4, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w135 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0010_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd5, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w136 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0010_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd6, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w137 = {1'b0, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0010_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'd7, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 13'h0002, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 2'b00, 1'b0, 4'b0000};
assign w138 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0010_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b00, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};
assign w139 = {1'b1, 1'b0, 1'b0, 8'h00, 5'b00011, 3'b000, 1'b0, 1'b0, 37'b0_0010_0000_0000_0000_0000_0000_0000_0000_0001, 18'b000000000_0_0_00_0_0_0_0_0, 2'b00, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, 2'b10, 3'b000, 3'b000, 3'b101, 3'b000, 3'b011, 3'b000, 3'b000, 3'b000, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 13'h0100, 13'h0001, 13'h0001, 13'h0001, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 2'b01, 2'b00, 2'b01, 1'b0, 4'b0000};

endmodule