module length_data(
    output wire [3071:0] out
);
    wire [7:0]wire0, wire1, wire2, wire3, wire4, wire5, wire6, wire7, wire8, wire9, wire10, wire11, wire12, wire13, wire14, wire15, wire16, wire17, wire18, wire19, wire20, wire21, wire22, wire23, wire24, wire25, wire26, wire27, wire28, wire29, wire30, wire31, wire32, wire33, wire34, wire35, wire36, wire37, wire38, wire39, wire40, wire41, wire42, wire43, wire44, wire45, wire46, wire47, wire48, wire49, wire50, wire51, wire52, wire53, wire54, wire55, wire56, wire57, wire58, wire59, wire60, wire61, wire62, wire63, wire64, wire65, wire66, wire67, wire68, wire69, wire70, wire71, wire72, wire73, wire74, wire75, wire76, wire77, wire78, wire79, wire80, wire81, wire82, wire83, wire84, wire85, wire86, wire87, wire88, wire89, wire90, wire91, wire92, wire93, wire94, wire95, wire96, wire97, wire98, wire99, wire100, wire101, wire102, wire103, wire104, wire105, wire106, wire107, wire108, wire109, wire110, wire111, wire112, wire113, wire114, wire115, wire116, wire117, wire118, wire119, wire120, wire121, wire122, wire123, wire124, wire125, wire126, wire127, wire128, wire129, wire130, wire131, wire132, wire133, wire134, wire135, wire136, wire137, wire138, wire139, wire140, wire141, wire142, wire143, wire144, wire145, wire146, wire147, wire148, wire149, wire150, wire151, wire152, wire153, wire154, wire155, wire156, wire157, wire158, wire159, wire160, wire161, wire162, wire163, wire164, wire165, wire166, wire167, wire168, wire169, wire170, wire171, wire172, wire173, wire174, wire175, wire176, wire177, wire178, wire179, wire180, wire181, wire182, wire183, wire184, wire185, wire186, wire187, wire188, wire189, wire190, wire191, wire192, wire193, wire194, wire195, wire196, wire197, wire198, wire199, wire200, wire201, wire202, wire203, wire204, wire205, wire206, wire207, wire208, wire209, wire210, wire211, wire212, wire213, wire214, wire215, wire216, wire217, wire218, wire219, wire220, wire221, wire222, wire223, wire224, wire225, wire226, wire227, wire228, wire229, wire230, wire231, wire232, wire233, wire234, wire235, wire236, wire237, wire238, wire239, wire240, wire241, wire242, wire243, wire244, wire245, wire246, wire247, wire248, wire249, wire250, wire251, wire252, wire253, wire254, wire255, wire256, wire257, wire258, wire259, wire260, wire261, wire262, wire263, wire264, wire265, wire266, wire267, wire268, wire269, wire270, wire271, wire272, wire273, wire274, wire275, wire276, wire277, wire278, wire279, wire280, wire281, wire282, wire283, wire284, wire285, wire286, wire287, wire288, wire289, wire290, wire291, wire292, wire293, wire294, wire295, wire296, wire297, wire298, wire299, wire300, wire301, wire302, wire303, wire304, wire305, wire306, wire307, wire308, wire309, wire310, wire311, wire312, wire313, wire314, wire315, wire316, wire317, wire318, wire319, wire320, wire321, wire322, wire323, wire324, wire325, wire326, wire327, wire328, wire329, wire330, wire331, wire332, wire333, wire334, wire335, wire336, wire337, wire338, wire339, wire340, wire341, wire342, wire343, wire344, wire345, wire346, wire347, wire348, wire349, wire350, wire351, wire352, wire353, wire354, wire355, wire356, wire357, wire358, wire359, wire360, wire361, wire362, wire363, wire364, wire365, wire366, wire367, wire368, wire369, wire370, wire371, wire372, wire373, wire374, wire375, wire376, wire377, wire378, wire379, wire380, wire381, wire382, wire383;
    assign wire0 = {8'd1};
    assign wire1 = {8'd2};
    assign wire2 = {8'd3};
    assign wire3 = {8'd4};
    assign wire4 = {8'd2};
    assign wire5 = {8'd3};
    assign wire6 = {8'd4};
    assign wire7 = {8'd5};
    assign wire8 = {8'd2};
    assign wire9 = {8'd3};
    assign wire10 = {8'd4};
    assign wire11 = {8'd5};
    assign wire12 = {8'd3};
    assign wire13 = {8'd4};
    assign wire14 = {8'd5};
    assign wire15 = {8'd6};
    assign wire16 = {8'd1};
    assign wire17 = {8'd2};
    assign wire18 = {8'd3};
    assign wire19 = {8'd4};
    assign wire20 = {8'd2};
    assign wire21 = {8'd3};
    assign wire22 = {8'd4};
    assign wire23 = {8'd5};
    assign wire24 = {8'd3};
    assign wire25 = {8'd4};
    assign wire26 = {8'd5};
    assign wire27 = {8'd6};
    assign wire28 = {8'd4};
    assign wire29 = {8'd5};
    assign wire30 = {8'd6};
    assign wire31 = {8'd7};
    assign wire32 = {8'd1};
    assign wire33 = {8'd2};
    assign wire34 = {8'd3};
    assign wire35 = {8'd4};
    assign wire36 = {8'd2};
    assign wire37 = {8'd3};
    assign wire38 = {8'd4};
    assign wire39 = {8'd5};
    assign wire40 = {8'd5};
    assign wire41 = {8'd6};
    assign wire42 = {8'd7};
    assign wire43 = {8'd8};
    assign wire44 = {8'd6};
    assign wire45 = {8'd7};
    assign wire46 = {8'd8};
    assign wire47 = {8'd9};
    assign wire48 = {8'd1};
    assign wire49 = {8'd2};
    assign wire50 = {8'd3};
    assign wire51 = {8'd4};
    assign wire52 = {8'd2};
    assign wire53 = {8'd3};
    assign wire54 = {8'd4};
    assign wire55 = {8'd5};
    assign wire56 = {8'd7};
    assign wire57 = {8'd8};
    assign wire58 = {8'd9};
    assign wire59 = {8'd10};
    assign wire60 = {8'd8};
    assign wire61 = {8'd9};
    assign wire62 = {8'd10};
    assign wire63 = {8'd11};
    assign wire64 = {8'd2};
    assign wire65 = {8'd3};
    assign wire66 = {8'd4};
    assign wire67 = {8'd5};
    assign wire68 = {8'd3};
    assign wire69 = {8'd4};
    assign wire70 = {8'd5};
    assign wire71 = {8'd6};
    assign wire72 = {8'd3};
    assign wire73 = {8'd4};
    assign wire74 = {8'd5};
    assign wire75 = {8'd6};
    assign wire76 = {8'd4};
    assign wire77 = {8'd5};
    assign wire78 = {8'd6};
    assign wire79 = {8'd7};
    assign wire80 = {8'd2};
    assign wire81 = {8'd3};
    assign wire82 = {8'd4};
    assign wire83 = {8'd5};
    assign wire84 = {8'd3};
    assign wire85 = {8'd4};
    assign wire86 = {8'd5};
    assign wire87 = {8'd6};
    assign wire88 = {8'd4};
    assign wire89 = {8'd5};
    assign wire90 = {8'd6};
    assign wire91 = {8'd7};
    assign wire92 = {8'd5};
    assign wire93 = {8'd6};
    assign wire94 = {8'd7};
    assign wire95 = {8'd8};
    assign wire96 = {8'd2};
    assign wire97 = {8'd3};
    assign wire98 = {8'd4};
    assign wire99 = {8'd5};
    assign wire100 = {8'd3};
    assign wire101 = {8'd4};
    assign wire102 = {8'd5};
    assign wire103 = {8'd6};
    assign wire104 = {8'd6};
    assign wire105 = {8'd7};
    assign wire106 = {8'd8};
    assign wire107 = {8'd9};
    assign wire108 = {8'd7};
    assign wire109 = {8'd8};
    assign wire110 = {8'd9};
    assign wire111 = {8'd10};
    assign wire112 = {8'd2};
    assign wire113 = {8'd3};
    assign wire114 = {8'd4};
    assign wire115 = {8'd5};
    assign wire116 = {8'd3};
    assign wire117 = {8'd4};
    assign wire118 = {8'd5};
    assign wire119 = {8'd6};
    assign wire120 = {8'd8};
    assign wire121 = {8'd9};
    assign wire122 = {8'd10};
    assign wire123 = {8'd11};
    assign wire124 = {8'd9};
    assign wire125 = {8'd10};
    assign wire126 = {8'd11};
    assign wire127 = {8'd12};
    assign wire128 = {8'd3};
    assign wire129 = {8'd4};
    assign wire130 = {8'd5};
    assign wire131 = {8'd6};
    assign wire132 = {8'd4};
    assign wire133 = {8'd5};
    assign wire134 = {8'd6};
    assign wire135 = {8'd7};
    assign wire136 = {8'd4};
    assign wire137 = {8'd5};
    assign wire138 = {8'd6};
    assign wire139 = {8'd7};
    assign wire140 = {8'd5};
    assign wire141 = {8'd6};
    assign wire142 = {8'd7};
    assign wire143 = {8'd8};
    assign wire144 = {8'd3};
    assign wire145 = {8'd4};
    assign wire146 = {8'd5};
    assign wire147 = {8'd6};
    assign wire148 = {8'd4};
    assign wire149 = {8'd5};
    assign wire150 = {8'd6};
    assign wire151 = {8'd7};
    assign wire152 = {8'd5};
    assign wire153 = {8'd6};
    assign wire154 = {8'd7};
    assign wire155 = {8'd8};
    assign wire156 = {8'd6};
    assign wire157 = {8'd7};
    assign wire158 = {8'd8};
    assign wire159 = {8'd9};
    assign wire160 = {8'd3};
    assign wire161 = {8'd4};
    assign wire162 = {8'd5};
    assign wire163 = {8'd6};
    assign wire164 = {8'd4};
    assign wire165 = {8'd5};
    assign wire166 = {8'd6};
    assign wire167 = {8'd7};
    assign wire168 = {8'd7};
    assign wire169 = {8'd8};
    assign wire170 = {8'd9};
    assign wire171 = {8'd10};
    assign wire172 = {8'd8};
    assign wire173 = {8'd9};
    assign wire174 = {8'd10};
    assign wire175 = {8'd11};
    assign wire176 = {8'd3};
    assign wire177 = {8'd4};
    assign wire178 = {8'd5};
    assign wire179 = {8'd6};
    assign wire180 = {8'd4};
    assign wire181 = {8'd5};
    assign wire182 = {8'd6};
    assign wire183 = {8'd7};
    assign wire184 = {8'd9};
    assign wire185 = {8'd10};
    assign wire186 = {8'd11};
    assign wire187 = {8'd12};
    assign wire188 = {8'd10};
    assign wire189 = {8'd11};
    assign wire190 = {8'd12};
    assign wire191 = {8'd13};
    assign wire192 = {8'd4};
    assign wire193 = {8'd5};
    assign wire194 = {8'd6};
    assign wire195 = {8'd7};
    assign wire196 = {8'd5};
    assign wire197 = {8'd6};
    assign wire198 = {8'd7};
    assign wire199 = {8'd8};
    assign wire200 = {8'd5};
    assign wire201 = {8'd6};
    assign wire202 = {8'd7};
    assign wire203 = {8'd8};
    assign wire204 = {8'd6};
    assign wire205 = {8'd7};
    assign wire206 = {8'd8};
    assign wire207 = {8'd9};
    assign wire208 = {8'd4};
    assign wire209 = {8'd5};
    assign wire210 = {8'd6};
    assign wire211 = {8'd7};
    assign wire212 = {8'd5};
    assign wire213 = {8'd6};
    assign wire214 = {8'd7};
    assign wire215 = {8'd8};
    assign wire216 = {8'd6};
    assign wire217 = {8'd7};
    assign wire218 = {8'd8};
    assign wire219 = {8'd9};
    assign wire220 = {8'd7};
    assign wire221 = {8'd8};
    assign wire222 = {8'd9};
    assign wire223 = {8'd10};
    assign wire224 = {8'd4};
    assign wire225 = {8'd5};
    assign wire226 = {8'd6};
    assign wire227 = {8'd7};
    assign wire228 = {8'd5};
    assign wire229 = {8'd6};
    assign wire230 = {8'd7};
    assign wire231 = {8'd8};
    assign wire232 = {8'd8};
    assign wire233 = {8'd9};
    assign wire234 = {8'd10};
    assign wire235 = {8'd11};
    assign wire236 = {8'd9};
    assign wire237 = {8'd10};
    assign wire238 = {8'd11};
    assign wire239 = {8'd12};
    assign wire240 = {8'd4};
    assign wire241 = {8'd5};
    assign wire242 = {8'd6};
    assign wire243 = {8'd7};
    assign wire244 = {8'd5};
    assign wire245 = {8'd6};
    assign wire246 = {8'd7};
    assign wire247 = {8'd8};
    assign wire248 = {8'd10};
    assign wire249 = {8'd11};
    assign wire250 = {8'd12};
    assign wire251 = {8'd13};
    assign wire252 = {8'd11};
    assign wire253 = {8'd12};
    assign wire254 = {8'd13};
    assign wire255 = {8'd14};
    assign wire256 = {8'd6};
    assign wire257 = {8'd7};
    assign wire258 = {8'd8};
    assign wire259 = {8'd9};
    assign wire260 = {8'd7};
    assign wire261 = {8'd8};
    assign wire262 = {8'd9};
    assign wire263 = {8'd10};
    assign wire264 = {8'd7};
    assign wire265 = {8'd8};
    assign wire266 = {8'd9};
    assign wire267 = {8'd10};
    assign wire268 = {8'd8};
    assign wire269 = {8'd9};
    assign wire270 = {8'd10};
    assign wire271 = {8'd11};
    assign wire272 = {8'd6};
    assign wire273 = {8'd7};
    assign wire274 = {8'd8};
    assign wire275 = {8'd9};
    assign wire276 = {8'd7};
    assign wire277 = {8'd8};
    assign wire278 = {8'd9};
    assign wire279 = {8'd10};
    assign wire280 = {8'd8};
    assign wire281 = {8'd9};
    assign wire282 = {8'd10};
    assign wire283 = {8'd11};
    assign wire284 = {8'd9};
    assign wire285 = {8'd10};
    assign wire286 = {8'd11};
    assign wire287 = {8'd12};
    assign wire288 = {8'd6};
    assign wire289 = {8'd7};
    assign wire290 = {8'd8};
    assign wire291 = {8'd9};
    assign wire292 = {8'd7};
    assign wire293 = {8'd8};
    assign wire294 = {8'd9};
    assign wire295 = {8'd10};
    assign wire296 = {8'd10};
    assign wire297 = {8'd11};
    assign wire298 = {8'd12};
    assign wire299 = {8'd13};
    assign wire300 = {8'd11};
    assign wire301 = {8'd12};
    assign wire302 = {8'd13};
    assign wire303 = {8'd14};
    assign wire304 = {8'd6};
    assign wire305 = {8'd7};
    assign wire306 = {8'd8};
    assign wire307 = {8'd9};
    assign wire308 = {8'd7};
    assign wire309 = {8'd8};
    assign wire310 = {8'd9};
    assign wire311 = {8'd10};
    assign wire312 = {8'd12};
    assign wire313 = {8'd13};
    assign wire314 = {8'd14};
    assign wire315 = {8'd15};
    assign wire316 = {8'd13};
    assign wire317 = {8'd14};
    assign wire318 = {8'd15};
    assign wire319 = {8'd16};
    assign wire320 = {8'd7};
    assign wire321 = {8'd8};
    assign wire322 = {8'd9};
    assign wire323 = {8'd10};
    assign wire324 = {8'd8};
    assign wire325 = {8'd9};
    assign wire326 = {8'd10};
    assign wire327 = {8'd11};
    assign wire328 = {8'd8};
    assign wire329 = {8'd9};
    assign wire330 = {8'd10};
    assign wire331 = {8'd11};
    assign wire332 = {8'd9};
    assign wire333 = {8'd10};
    assign wire334 = {8'd11};
    assign wire335 = {8'd12};
    assign wire336 = {8'd7};
    assign wire337 = {8'd8};
    assign wire338 = {8'd9};
    assign wire339 = {8'd10};
    assign wire340 = {8'd8};
    assign wire341 = {8'd9};
    assign wire342 = {8'd10};
    assign wire343 = {8'd11};
    assign wire344 = {8'd9};
    assign wire345 = {8'd10};
    assign wire346 = {8'd11};
    assign wire347 = {8'd12};
    assign wire348 = {8'd10};
    assign wire349 = {8'd11};
    assign wire350 = {8'd12};
    assign wire351 = {8'd13};
    assign wire352 = {8'd7};
    assign wire353 = {8'd8};
    assign wire354 = {8'd9};
    assign wire355 = {8'd10};
    assign wire356 = {8'd8};
    assign wire357 = {8'd9};
    assign wire358 = {8'd10};
    assign wire359 = {8'd11};
    assign wire360 = {8'd11};
    assign wire361 = {8'd12};
    assign wire362 = {8'd13};
    assign wire363 = {8'd14};
    assign wire364 = {8'd12};
    assign wire365 = {8'd13};
    assign wire366 = {8'd14};
    assign wire367 = {8'd15};
    assign wire368 = {8'd7};
    assign wire369 = {8'd8};
    assign wire370 = {8'd9};
    assign wire371 = {8'd10};
    assign wire372 = {8'd8};
    assign wire373 = {8'd9};
    assign wire374 = {8'd10};
    assign wire375 = {8'd11};
    assign wire376 = {8'd13};
    assign wire377 = {8'd14};
    assign wire378 = {8'd15};
    assign wire379 = {8'd16};
    assign wire380 = {8'd14};
    assign wire381 = {8'd15};
    assign wire382 = {8'd16};
    assign wire383 = {8'd17};
    wire [3071:0] data_concat;
    assign data_concat = {wire383, wire382, wire381, wire380, wire379, wire378, wire377, wire376, wire375, wire374, wire373, wire372, wire371, wire370, wire369, wire368, wire367, wire366, wire365, wire364, wire363, wire362, wire361, wire360, wire359, wire358, wire357, wire356, wire355, wire354, wire353, wire352, wire351, wire350, wire349, wire348, wire347, wire346, wire345, wire344, wire343, wire342, wire341, wire340, wire339, wire338, wire337, wire336, wire335, wire334, wire333, wire332, wire331, wire330, wire329, wire328, wire327, wire326, wire325, wire324, wire323, wire322, wire321, wire320, wire319, wire318, wire317, wire316, wire315, wire314, wire313, wire312, wire311, wire310, wire309, wire308, wire307, wire306, wire305, wire304, wire303, wire302, wire301, wire300, wire299, wire298, wire297, wire296, wire295, wire294, wire293, wire292, wire291, wire290, wire289, wire288, wire287, wire286, wire285, wire284, wire283, wire282, wire281, wire280, wire279, wire278, wire277, wire276, wire275, wire274, wire273, wire272, wire271, wire270, wire269, wire268, wire267, wire266, wire265, wire264, wire263, wire262, wire261, wire260, wire259, wire258, wire257, wire256, wire255, wire254, wire253, wire252, wire251, wire250, wire249, wire248, wire247, wire246, wire245, wire244, wire243, wire242, wire241, wire240, wire239, wire238, wire237, wire236, wire235, wire234, wire233, wire232, wire231, wire230, wire229, wire228, wire227, wire226, wire225, wire224, wire223, wire222, wire221, wire220, wire219, wire218, wire217, wire216, wire215, wire214, wire213, wire212, wire211, wire210, wire209, wire208, wire207, wire206, wire205, wire204, wire203, wire202, wire201, wire200, wire199, wire198, wire197, wire196, wire195, wire194, wire193, wire192, wire191, wire190, wire189, wire188, wire187, wire186, wire185, wire184, wire183, wire182, wire181, wire180, wire179, wire178, wire177, wire176, wire175, wire174, wire173, wire172, wire171, wire170, wire169, wire168, wire167, wire166, wire165, wire164, wire163, wire162, wire161, wire160, wire159, wire158, wire157, wire156, wire155, wire154, wire153, wire152, wire151, wire150, wire149, wire148, wire147, wire146, wire145, wire144, wire143, wire142, wire141, wire140, wire139, wire138, wire137, wire136, wire135, wire134, wire133, wire132, wire131, wire130, wire129, wire128, wire127, wire126, wire125, wire124, wire123, wire122, wire121, wire120, wire119, wire118, wire117, wire116, wire115, wire114, wire113, wire112, wire111, wire110, wire109, wire108, wire107, wire106, wire105, wire104, wire103, wire102, wire101, wire100, wire99, wire98, wire97, wire96, wire95, wire94, wire93, wire92, wire91, wire90, wire89, wire88, wire87, wire86, wire85, wire84, wire83, wire82, wire81, wire80, wire79, wire78, wire77, wire76, wire75, wire74, wire73, wire72, wire71, wire70, wire69, wire68, wire67, wire66, wire65, wire64, wire63, wire62, wire61, wire60, wire59, wire58, wire57, wire56, wire55, wire54, wire53, wire52, wire51, wire50, wire49, wire48, wire47, wire46, wire45, wire44, wire43, wire42, wire41, wire40, wire39, wire38, wire37, wire36, wire35, wire34, wire33, wire32, wire31, wire30, wire29, wire28, wire27, wire26, wire25, wire24, wire23, wire22, wire21, wire20, wire19, wire18, wire17, wire16, wire15, wire14, wire13, wire12, wire11, wire10, wire9, wire8, wire7, wire6, wire5, wire4, wire3, wire2, wire1, wire0};
    assign out = data_concat;


endmodule

