module length_data(
    output wire [40959:0] out
);
    wire [9:0] wire0, wire1, wire2, wire3, wire4, wire5, wire6, wire7, wire8, wire9, wire10, wire11, wire12, wire13, wire14, wire15, wire16, wire17, wire18, wire19, wire20, wire21, wire22, wire23, wire24, wire25, wire26, wire27, wire28, wire29, wire30, wire31, wire32, wire33, wire34, wire35, wire36, wire37, wire38, wire39, wire40, wire41, wire42, wire43, wire44, wire45, wire46, wire47, wire48, wire49, wire50, wire51, wire52, wire53, wire54, wire55, wire56, wire57, wire58, wire59, wire60, wire61, wire62, wire63, wire64, wire65, wire66, wire67, wire68, wire69, wire70, wire71, wire72, wire73, wire74, wire75, wire76, wire77, wire78, wire79, wire80, wire81, wire82, wire83, wire84, wire85, wire86, wire87, wire88, wire89, wire90, wire91, wire92, wire93, wire94, wire95, wire96, wire97, wire98, wire99, wire100, wire101, wire102, wire103, wire104, wire105, wire106, wire107, wire108, wire109, wire110, wire111, wire112, wire113, wire114, wire115, wire116, wire117, wire118, wire119, wire120, wire121, wire122, wire123, wire124, wire125, wire126, wire127, wire128, wire129, wire130, wire131, wire132, wire133, wire134, wire135, wire136, wire137, wire138, wire139, wire140, wire141, wire142, wire143, wire144, wire145, wire146, wire147, wire148, wire149, wire150, wire151, wire152, wire153, wire154, wire155, wire156, wire157, wire158, wire159, wire160, wire161, wire162, wire163, wire164, wire165, wire166, wire167, wire168, wire169, wire170, wire171, wire172, wire173, wire174, wire175, wire176, wire177, wire178, wire179, wire180, wire181, wire182, wire183, wire184, wire185, wire186, wire187, wire188, wire189, wire190, wire191, wire192, wire193, wire194, wire195, wire196, wire197, wire198, wire199, wire200, wire201, wire202, wire203, wire204, wire205, wire206, wire207, wire208, wire209, wire210, wire211, wire212, wire213, wire214, wire215, wire216, wire217, wire218, wire219, wire220, wire221, wire222, wire223, wire224, wire225, wire226, wire227, wire228, wire229, wire230, wire231, wire232, wire233, wire234, wire235, wire236, wire237, wire238, wire239, wire240, wire241, wire242, wire243, wire244, wire245, wire246, wire247, wire248, wire249, wire250, wire251, wire252, wire253, wire254, wire255, wire256, wire257, wire258, wire259, wire260, wire261, wire262, wire263, wire264, wire265, wire266, wire267, wire268, wire269, wire270, wire271, wire272, wire273, wire274, wire275, wire276, wire277, wire278, wire279, wire280, wire281, wire282, wire283, wire284, wire285, wire286, wire287, wire288, wire289, wire290, wire291, wire292, wire293, wire294, wire295, wire296, wire297, wire298, wire299, wire300, wire301, wire302, wire303, wire304, wire305, wire306, wire307, wire308, wire309, wire310, wire311, wire312, wire313, wire314, wire315, wire316, wire317, wire318, wire319, wire320, wire321, wire322, wire323, wire324, wire325, wire326, wire327, wire328, wire329, wire330, wire331, wire332, wire333, wire334, wire335, wire336, wire337, wire338, wire339, wire340, wire341, wire342, wire343, wire344, wire345, wire346, wire347, wire348, wire349, wire350, wire351, wire352, wire353, wire354, wire355, wire356, wire357, wire358, wire359, wire360, wire361, wire362, wire363, wire364, wire365, wire366, wire367, wire368, wire369, wire370, wire371, wire372, wire373, wire374, wire375, wire376, wire377, wire378, wire379, wire380, wire381, wire382, wire383, wire384, wire385, wire386, wire387, wire388, wire389, wire390, wire391, wire392, wire393, wire394, wire395, wire396, wire397, wire398, wire399, wire400, wire401, wire402, wire403, wire404, wire405, wire406, wire407, wire408, wire409, wire410, wire411, wire412, wire413, wire414, wire415, wire416, wire417, wire418, wire419, wire420, wire421, wire422, wire423, wire424, wire425, wire426, wire427, wire428, wire429, wire430, wire431, wire432, wire433, wire434, wire435, wire436, wire437, wire438, wire439, wire440, wire441, wire442, wire443, wire444, wire445, wire446, wire447, wire448, wire449, wire450, wire451, wire452, wire453, wire454, wire455, wire456, wire457, wire458, wire459, wire460, wire461, wire462, wire463, wire464, wire465, wire466, wire467, wire468, wire469, wire470, wire471, wire472, wire473, wire474, wire475, wire476, wire477, wire478, wire479, wire480, wire481, wire482, wire483, wire484, wire485, wire486, wire487, wire488, wire489, wire490, wire491, wire492, wire493, wire494, wire495, wire496, wire497, wire498, wire499, wire500, wire501, wire502, wire503, wire504, wire505, wire506, wire507, wire508, wire509, wire510, wire511, wire512, wire513, wire514, wire515, wire516, wire517, wire518, wire519, wire520, wire521, wire522, wire523, wire524, wire525, wire526, wire527, wire528, wire529, wire530, wire531, wire532, wire533, wire534, wire535, wire536, wire537, wire538, wire539, wire540, wire541, wire542, wire543, wire544, wire545, wire546, wire547, wire548, wire549, wire550, wire551, wire552, wire553, wire554, wire555, wire556, wire557, wire558, wire559, wire560, wire561, wire562, wire563, wire564, wire565, wire566, wire567, wire568, wire569, wire570, wire571, wire572, wire573, wire574, wire575, wire576, wire577, wire578, wire579, wire580, wire581, wire582, wire583, wire584, wire585, wire586, wire587, wire588, wire589, wire590, wire591, wire592, wire593, wire594, wire595, wire596, wire597, wire598, wire599, wire600, wire601, wire602, wire603, wire604, wire605, wire606, wire607, wire608, wire609, wire610, wire611, wire612, wire613, wire614, wire615, wire616, wire617, wire618, wire619, wire620, wire621, wire622, wire623, wire624, wire625, wire626, wire627, wire628, wire629, wire630, wire631, wire632, wire633, wire634, wire635, wire636, wire637, wire638, wire639, wire640, wire641, wire642, wire643, wire644, wire645, wire646, wire647, wire648, wire649, wire650, wire651, wire652, wire653, wire654, wire655, wire656, wire657, wire658, wire659, wire660, wire661, wire662, wire663, wire664, wire665, wire666, wire667, wire668, wire669, wire670, wire671, wire672, wire673, wire674, wire675, wire676, wire677, wire678, wire679, wire680, wire681, wire682, wire683, wire684, wire685, wire686, wire687, wire688, wire689, wire690, wire691, wire692, wire693, wire694, wire695, wire696, wire697, wire698, wire699, wire700, wire701, wire702, wire703, wire704, wire705, wire706, wire707, wire708, wire709, wire710, wire711, wire712, wire713, wire714, wire715, wire716, wire717, wire718, wire719, wire720, wire721, wire722, wire723, wire724, wire725, wire726, wire727, wire728, wire729, wire730, wire731, wire732, wire733, wire734, wire735, wire736, wire737, wire738, wire739, wire740, wire741, wire742, wire743, wire744, wire745, wire746, wire747, wire748, wire749, wire750, wire751, wire752, wire753, wire754, wire755, wire756, wire757, wire758, wire759, wire760, wire761, wire762, wire763, wire764, wire765, wire766, wire767, wire768, wire769, wire770, wire771, wire772, wire773, wire774, wire775, wire776, wire777, wire778, wire779, wire780, wire781, wire782, wire783, wire784, wire785, wire786, wire787, wire788, wire789, wire790, wire791, wire792, wire793, wire794, wire795, wire796, wire797, wire798, wire799, wire800, wire801, wire802, wire803, wire804, wire805, wire806, wire807, wire808, wire809, wire810, wire811, wire812, wire813, wire814, wire815, wire816, wire817, wire818, wire819, wire820, wire821, wire822, wire823, wire824, wire825, wire826, wire827, wire828, wire829, wire830, wire831, wire832, wire833, wire834, wire835, wire836, wire837, wire838, wire839, wire840, wire841, wire842, wire843, wire844, wire845, wire846, wire847, wire848, wire849, wire850, wire851, wire852, wire853, wire854, wire855, wire856, wire857, wire858, wire859, wire860, wire861, wire862, wire863, wire864, wire865, wire866, wire867, wire868, wire869, wire870, wire871, wire872, wire873, wire874, wire875, wire876, wire877, wire878, wire879, wire880, wire881, wire882, wire883, wire884, wire885, wire886, wire887, wire888, wire889, wire890, wire891, wire892, wire893, wire894, wire895, wire896, wire897, wire898, wire899, wire900, wire901, wire902, wire903, wire904, wire905, wire906, wire907, wire908, wire909, wire910, wire911, wire912, wire913, wire914, wire915, wire916, wire917, wire918, wire919, wire920, wire921, wire922, wire923, wire924, wire925, wire926, wire927, wire928, wire929, wire930, wire931, wire932, wire933, wire934, wire935, wire936, wire937, wire938, wire939, wire940, wire941, wire942, wire943, wire944, wire945, wire946, wire947, wire948, wire949, wire950, wire951, wire952, wire953, wire954, wire955, wire956, wire957, wire958, wire959, wire960, wire961, wire962, wire963, wire964, wire965, wire966, wire967, wire968, wire969, wire970, wire971, wire972, wire973, wire974, wire975, wire976, wire977, wire978, wire979, wire980, wire981, wire982, wire983, wire984, wire985, wire986, wire987, wire988, wire989, wire990, wire991, wire992, wire993, wire994, wire995, wire996, wire997, wire998, wire999, wire1000, wire1001, wire1002, wire1003, wire1004, wire1005, wire1006, wire1007, wire1008, wire1009, wire1010, wire1011, wire1012, wire1013, wire1014, wire1015, wire1016, wire1017, wire1018, wire1019, wire1020, wire1021, wire1022, wire1023, wire1024, wire1025, wire1026, wire1027, wire1028, wire1029, wire1030, wire1031, wire1032, wire1033, wire1034, wire1035, wire1036, wire1037, wire1038, wire1039, wire1040, wire1041, wire1042, wire1043, wire1044, wire1045, wire1046, wire1047, wire1048, wire1049, wire1050, wire1051, wire1052, wire1053, wire1054, wire1055, wire1056, wire1057, wire1058, wire1059, wire1060, wire1061, wire1062, wire1063, wire1064, wire1065, wire1066, wire1067, wire1068, wire1069, wire1070, wire1071, wire1072, wire1073, wire1074, wire1075, wire1076, wire1077, wire1078, wire1079, wire1080, wire1081, wire1082, wire1083, wire1084, wire1085, wire1086, wire1087, wire1088, wire1089, wire1090, wire1091, wire1092, wire1093, wire1094, wire1095, wire1096, wire1097, wire1098, wire1099, wire1100, wire1101, wire1102, wire1103, wire1104, wire1105, wire1106, wire1107, wire1108, wire1109, wire1110, wire1111, wire1112, wire1113, wire1114, wire1115, wire1116, wire1117, wire1118, wire1119, wire1120, wire1121, wire1122, wire1123, wire1124, wire1125, wire1126, wire1127, wire1128, wire1129, wire1130, wire1131, wire1132, wire1133, wire1134, wire1135, wire1136, wire1137, wire1138, wire1139, wire1140, wire1141, wire1142, wire1143, wire1144, wire1145, wire1146, wire1147, wire1148, wire1149, wire1150, wire1151, wire1152, wire1153, wire1154, wire1155, wire1156, wire1157, wire1158, wire1159, wire1160, wire1161, wire1162, wire1163, wire1164, wire1165, wire1166, wire1167, wire1168, wire1169, wire1170, wire1171, wire1172, wire1173, wire1174, wire1175, wire1176, wire1177, wire1178, wire1179, wire1180, wire1181, wire1182, wire1183, wire1184, wire1185, wire1186, wire1187, wire1188, wire1189, wire1190, wire1191, wire1192, wire1193, wire1194, wire1195, wire1196, wire1197, wire1198, wire1199, wire1200, wire1201, wire1202, wire1203, wire1204, wire1205, wire1206, wire1207, wire1208, wire1209, wire1210, wire1211, wire1212, wire1213, wire1214, wire1215, wire1216, wire1217, wire1218, wire1219, wire1220, wire1221, wire1222, wire1223, wire1224, wire1225, wire1226, wire1227, wire1228, wire1229, wire1230, wire1231, wire1232, wire1233, wire1234, wire1235, wire1236, wire1237, wire1238, wire1239, wire1240, wire1241, wire1242, wire1243, wire1244, wire1245, wire1246, wire1247, wire1248, wire1249, wire1250, wire1251, wire1252, wire1253, wire1254, wire1255, wire1256, wire1257, wire1258, wire1259, wire1260, wire1261, wire1262, wire1263, wire1264, wire1265, wire1266, wire1267, wire1268, wire1269, wire1270, wire1271, wire1272, wire1273, wire1274, wire1275, wire1276, wire1277, wire1278, wire1279, wire1280, wire1281, wire1282, wire1283, wire1284, wire1285, wire1286, wire1287, wire1288, wire1289, wire1290, wire1291, wire1292, wire1293, wire1294, wire1295, wire1296, wire1297, wire1298, wire1299, wire1300, wire1301, wire1302, wire1303, wire1304, wire1305, wire1306, wire1307, wire1308, wire1309, wire1310, wire1311, wire1312, wire1313, wire1314, wire1315, wire1316, wire1317, wire1318, wire1319, wire1320, wire1321, wire1322, wire1323, wire1324, wire1325, wire1326, wire1327, wire1328, wire1329, wire1330, wire1331, wire1332, wire1333, wire1334, wire1335, wire1336, wire1337, wire1338, wire1339, wire1340, wire1341, wire1342, wire1343, wire1344, wire1345, wire1346, wire1347, wire1348, wire1349, wire1350, wire1351, wire1352, wire1353, wire1354, wire1355, wire1356, wire1357, wire1358, wire1359, wire1360, wire1361, wire1362, wire1363, wire1364, wire1365, wire1366, wire1367, wire1368, wire1369, wire1370, wire1371, wire1372, wire1373, wire1374, wire1375, wire1376, wire1377, wire1378, wire1379, wire1380, wire1381, wire1382, wire1383, wire1384, wire1385, wire1386, wire1387, wire1388, wire1389, wire1390, wire1391, wire1392, wire1393, wire1394, wire1395, wire1396, wire1397, wire1398, wire1399, wire1400, wire1401, wire1402, wire1403, wire1404, wire1405, wire1406, wire1407, wire1408, wire1409, wire1410, wire1411, wire1412, wire1413, wire1414, wire1415, wire1416, wire1417, wire1418, wire1419, wire1420, wire1421, wire1422, wire1423, wire1424, wire1425, wire1426, wire1427, wire1428, wire1429, wire1430, wire1431, wire1432, wire1433, wire1434, wire1435, wire1436, wire1437, wire1438, wire1439, wire1440, wire1441, wire1442, wire1443, wire1444, wire1445, wire1446, wire1447, wire1448, wire1449, wire1450, wire1451, wire1452, wire1453, wire1454, wire1455, wire1456, wire1457, wire1458, wire1459, wire1460, wire1461, wire1462, wire1463, wire1464, wire1465, wire1466, wire1467, wire1468, wire1469, wire1470, wire1471, wire1472, wire1473, wire1474, wire1475, wire1476, wire1477, wire1478, wire1479, wire1480, wire1481, wire1482, wire1483, wire1484, wire1485, wire1486, wire1487, wire1488, wire1489, wire1490, wire1491, wire1492, wire1493, wire1494, wire1495, wire1496, wire1497, wire1498, wire1499, wire1500, wire1501, wire1502, wire1503, wire1504, wire1505, wire1506, wire1507, wire1508, wire1509, wire1510, wire1511, wire1512, wire1513, wire1514, wire1515, wire1516, wire1517, wire1518, wire1519, wire1520, wire1521, wire1522, wire1523, wire1524, wire1525, wire1526, wire1527, wire1528, wire1529, wire1530, wire1531, wire1532, wire1533, wire1534, wire1535, wire1536, wire1537, wire1538, wire1539, wire1540, wire1541, wire1542, wire1543, wire1544, wire1545, wire1546, wire1547, wire1548, wire1549, wire1550, wire1551, wire1552, wire1553, wire1554, wire1555, wire1556, wire1557, wire1558, wire1559, wire1560, wire1561, wire1562, wire1563, wire1564, wire1565, wire1566, wire1567, wire1568, wire1569, wire1570, wire1571, wire1572, wire1573, wire1574, wire1575, wire1576, wire1577, wire1578, wire1579, wire1580, wire1581, wire1582, wire1583, wire1584, wire1585, wire1586, wire1587, wire1588, wire1589, wire1590, wire1591, wire1592, wire1593, wire1594, wire1595, wire1596, wire1597, wire1598, wire1599, wire1600, wire1601, wire1602, wire1603, wire1604, wire1605, wire1606, wire1607, wire1608, wire1609, wire1610, wire1611, wire1612, wire1613, wire1614, wire1615, wire1616, wire1617, wire1618, wire1619, wire1620, wire1621, wire1622, wire1623, wire1624, wire1625, wire1626, wire1627, wire1628, wire1629, wire1630, wire1631, wire1632, wire1633, wire1634, wire1635, wire1636, wire1637, wire1638, wire1639, wire1640, wire1641, wire1642, wire1643, wire1644, wire1645, wire1646, wire1647, wire1648, wire1649, wire1650, wire1651, wire1652, wire1653, wire1654, wire1655, wire1656, wire1657, wire1658, wire1659, wire1660, wire1661, wire1662, wire1663, wire1664, wire1665, wire1666, wire1667, wire1668, wire1669, wire1670, wire1671, wire1672, wire1673, wire1674, wire1675, wire1676, wire1677, wire1678, wire1679, wire1680, wire1681, wire1682, wire1683, wire1684, wire1685, wire1686, wire1687, wire1688, wire1689, wire1690, wire1691, wire1692, wire1693, wire1694, wire1695, wire1696, wire1697, wire1698, wire1699, wire1700, wire1701, wire1702, wire1703, wire1704, wire1705, wire1706, wire1707, wire1708, wire1709, wire1710, wire1711, wire1712, wire1713, wire1714, wire1715, wire1716, wire1717, wire1718, wire1719, wire1720, wire1721, wire1722, wire1723, wire1724, wire1725, wire1726, wire1727, wire1728, wire1729, wire1730, wire1731, wire1732, wire1733, wire1734, wire1735, wire1736, wire1737, wire1738, wire1739, wire1740, wire1741, wire1742, wire1743, wire1744, wire1745, wire1746, wire1747, wire1748, wire1749, wire1750, wire1751, wire1752, wire1753, wire1754, wire1755, wire1756, wire1757, wire1758, wire1759, wire1760, wire1761, wire1762, wire1763, wire1764, wire1765, wire1766, wire1767, wire1768, wire1769, wire1770, wire1771, wire1772, wire1773, wire1774, wire1775, wire1776, wire1777, wire1778, wire1779, wire1780, wire1781, wire1782, wire1783, wire1784, wire1785, wire1786, wire1787, wire1788, wire1789, wire1790, wire1791, wire1792, wire1793, wire1794, wire1795, wire1796, wire1797, wire1798, wire1799, wire1800, wire1801, wire1802, wire1803, wire1804, wire1805, wire1806, wire1807, wire1808, wire1809, wire1810, wire1811, wire1812, wire1813, wire1814, wire1815, wire1816, wire1817, wire1818, wire1819, wire1820, wire1821, wire1822, wire1823, wire1824, wire1825, wire1826, wire1827, wire1828, wire1829, wire1830, wire1831, wire1832, wire1833, wire1834, wire1835, wire1836, wire1837, wire1838, wire1839, wire1840, wire1841, wire1842, wire1843, wire1844, wire1845, wire1846, wire1847, wire1848, wire1849, wire1850, wire1851, wire1852, wire1853, wire1854, wire1855, wire1856, wire1857, wire1858, wire1859, wire1860, wire1861, wire1862, wire1863, wire1864, wire1865, wire1866, wire1867, wire1868, wire1869, wire1870, wire1871, wire1872, wire1873, wire1874, wire1875, wire1876, wire1877, wire1878, wire1879, wire1880, wire1881, wire1882, wire1883, wire1884, wire1885, wire1886, wire1887, wire1888, wire1889, wire1890, wire1891, wire1892, wire1893, wire1894, wire1895, wire1896, wire1897, wire1898, wire1899, wire1900, wire1901, wire1902, wire1903, wire1904, wire1905, wire1906, wire1907, wire1908, wire1909, wire1910, wire1911, wire1912, wire1913, wire1914, wire1915, wire1916, wire1917, wire1918, wire1919, wire1920, wire1921, wire1922, wire1923, wire1924, wire1925, wire1926, wire1927, wire1928, wire1929, wire1930, wire1931, wire1932, wire1933, wire1934, wire1935, wire1936, wire1937, wire1938, wire1939, wire1940, wire1941, wire1942, wire1943, wire1944, wire1945, wire1946, wire1947, wire1948, wire1949, wire1950, wire1951, wire1952, wire1953, wire1954, wire1955, wire1956, wire1957, wire1958, wire1959, wire1960, wire1961, wire1962, wire1963, wire1964, wire1965, wire1966, wire1967, wire1968, wire1969, wire1970, wire1971, wire1972, wire1973, wire1974, wire1975, wire1976, wire1977, wire1978, wire1979, wire1980, wire1981, wire1982, wire1983, wire1984, wire1985, wire1986, wire1987, wire1988, wire1989, wire1990, wire1991, wire1992, wire1993, wire1994, wire1995, wire1996, wire1997, wire1998, wire1999, wire2000, wire2001, wire2002, wire2003, wire2004, wire2005, wire2006, wire2007, wire2008, wire2009, wire2010, wire2011, wire2012, wire2013, wire2014, wire2015, wire2016, wire2017, wire2018, wire2019, wire2020, wire2021, wire2022, wire2023, wire2024, wire2025, wire2026, wire2027, wire2028, wire2029, wire2030, wire2031, wire2032, wire2033, wire2034, wire2035, wire2036, wire2037, wire2038, wire2039, wire2040, wire2041, wire2042, wire2043, wire2044, wire2045, wire2046, wire2047, wire2048, wire2049, wire2050, wire2051, wire2052, wire2053, wire2054, wire2055, wire2056, wire2057, wire2058, wire2059, wire2060, wire2061, wire2062, wire2063, wire2064, wire2065, wire2066, wire2067, wire2068, wire2069, wire2070, wire2071, wire2072, wire2073, wire2074, wire2075, wire2076, wire2077, wire2078, wire2079, wire2080, wire2081, wire2082, wire2083, wire2084, wire2085, wire2086, wire2087, wire2088, wire2089, wire2090, wire2091, wire2092, wire2093, wire2094, wire2095, wire2096, wire2097, wire2098, wire2099, wire2100, wire2101, wire2102, wire2103, wire2104, wire2105, wire2106, wire2107, wire2108, wire2109, wire2110, wire2111, wire2112, wire2113, wire2114, wire2115, wire2116, wire2117, wire2118, wire2119, wire2120, wire2121, wire2122, wire2123, wire2124, wire2125, wire2126, wire2127, wire2128, wire2129, wire2130, wire2131, wire2132, wire2133, wire2134, wire2135, wire2136, wire2137, wire2138, wire2139, wire2140, wire2141, wire2142, wire2143, wire2144, wire2145, wire2146, wire2147, wire2148, wire2149, wire2150, wire2151, wire2152, wire2153, wire2154, wire2155, wire2156, wire2157, wire2158, wire2159, wire2160, wire2161, wire2162, wire2163, wire2164, wire2165, wire2166, wire2167, wire2168, wire2169, wire2170, wire2171, wire2172, wire2173, wire2174, wire2175, wire2176, wire2177, wire2178, wire2179, wire2180, wire2181, wire2182, wire2183, wire2184, wire2185, wire2186, wire2187, wire2188, wire2189, wire2190, wire2191, wire2192, wire2193, wire2194, wire2195, wire2196, wire2197, wire2198, wire2199, wire2200, wire2201, wire2202, wire2203, wire2204, wire2205, wire2206, wire2207, wire2208, wire2209, wire2210, wire2211, wire2212, wire2213, wire2214, wire2215, wire2216, wire2217, wire2218, wire2219, wire2220, wire2221, wire2222, wire2223, wire2224, wire2225, wire2226, wire2227, wire2228, wire2229, wire2230, wire2231, wire2232, wire2233, wire2234, wire2235, wire2236, wire2237, wire2238, wire2239, wire2240, wire2241, wire2242, wire2243, wire2244, wire2245, wire2246, wire2247, wire2248, wire2249, wire2250, wire2251, wire2252, wire2253, wire2254, wire2255, wire2256, wire2257, wire2258, wire2259, wire2260, wire2261, wire2262, wire2263, wire2264, wire2265, wire2266, wire2267, wire2268, wire2269, wire2270, wire2271, wire2272, wire2273, wire2274, wire2275, wire2276, wire2277, wire2278, wire2279, wire2280, wire2281, wire2282, wire2283, wire2284, wire2285, wire2286, wire2287, wire2288, wire2289, wire2290, wire2291, wire2292, wire2293, wire2294, wire2295, wire2296, wire2297, wire2298, wire2299, wire2300, wire2301, wire2302, wire2303, wire2304, wire2305, wire2306, wire2307, wire2308, wire2309, wire2310, wire2311, wire2312, wire2313, wire2314, wire2315, wire2316, wire2317, wire2318, wire2319, wire2320, wire2321, wire2322, wire2323, wire2324, wire2325, wire2326, wire2327, wire2328, wire2329, wire2330, wire2331, wire2332, wire2333, wire2334, wire2335, wire2336, wire2337, wire2338, wire2339, wire2340, wire2341, wire2342, wire2343, wire2344, wire2345, wire2346, wire2347, wire2348, wire2349, wire2350, wire2351, wire2352, wire2353, wire2354, wire2355, wire2356, wire2357, wire2358, wire2359, wire2360, wire2361, wire2362, wire2363, wire2364, wire2365, wire2366, wire2367, wire2368, wire2369, wire2370, wire2371, wire2372, wire2373, wire2374, wire2375, wire2376, wire2377, wire2378, wire2379, wire2380, wire2381, wire2382, wire2383, wire2384, wire2385, wire2386, wire2387, wire2388, wire2389, wire2390, wire2391, wire2392, wire2393, wire2394, wire2395, wire2396, wire2397, wire2398, wire2399, wire2400, wire2401, wire2402, wire2403, wire2404, wire2405, wire2406, wire2407, wire2408, wire2409, wire2410, wire2411, wire2412, wire2413, wire2414, wire2415, wire2416, wire2417, wire2418, wire2419, wire2420, wire2421, wire2422, wire2423, wire2424, wire2425, wire2426, wire2427, wire2428, wire2429, wire2430, wire2431, wire2432, wire2433, wire2434, wire2435, wire2436, wire2437, wire2438, wire2439, wire2440, wire2441, wire2442, wire2443, wire2444, wire2445, wire2446, wire2447, wire2448, wire2449, wire2450, wire2451, wire2452, wire2453, wire2454, wire2455, wire2456, wire2457, wire2458, wire2459, wire2460, wire2461, wire2462, wire2463, wire2464, wire2465, wire2466, wire2467, wire2468, wire2469, wire2470, wire2471, wire2472, wire2473, wire2474, wire2475, wire2476, wire2477, wire2478, wire2479, wire2480, wire2481, wire2482, wire2483, wire2484, wire2485, wire2486, wire2487, wire2488, wire2489, wire2490, wire2491, wire2492, wire2493, wire2494, wire2495, wire2496, wire2497, wire2498, wire2499, wire2500, wire2501, wire2502, wire2503, wire2504, wire2505, wire2506, wire2507, wire2508, wire2509, wire2510, wire2511, wire2512, wire2513, wire2514, wire2515, wire2516, wire2517, wire2518, wire2519, wire2520, wire2521, wire2522, wire2523, wire2524, wire2525, wire2526, wire2527, wire2528, wire2529, wire2530, wire2531, wire2532, wire2533, wire2534, wire2535, wire2536, wire2537, wire2538, wire2539, wire2540, wire2541, wire2542, wire2543, wire2544, wire2545, wire2546, wire2547, wire2548, wire2549, wire2550, wire2551, wire2552, wire2553, wire2554, wire2555, wire2556, wire2557, wire2558, wire2559, wire2560, wire2561, wire2562, wire2563, wire2564, wire2565, wire2566, wire2567, wire2568, wire2569, wire2570, wire2571, wire2572, wire2573, wire2574, wire2575, wire2576, wire2577, wire2578, wire2579, wire2580, wire2581, wire2582, wire2583, wire2584, wire2585, wire2586, wire2587, wire2588, wire2589, wire2590, wire2591, wire2592, wire2593, wire2594, wire2595, wire2596, wire2597, wire2598, wire2599, wire2600, wire2601, wire2602, wire2603, wire2604, wire2605, wire2606, wire2607, wire2608, wire2609, wire2610, wire2611, wire2612, wire2613, wire2614, wire2615, wire2616, wire2617, wire2618, wire2619, wire2620, wire2621, wire2622, wire2623, wire2624, wire2625, wire2626, wire2627, wire2628, wire2629, wire2630, wire2631, wire2632, wire2633, wire2634, wire2635, wire2636, wire2637, wire2638, wire2639, wire2640, wire2641, wire2642, wire2643, wire2644, wire2645, wire2646, wire2647, wire2648, wire2649, wire2650, wire2651, wire2652, wire2653, wire2654, wire2655, wire2656, wire2657, wire2658, wire2659, wire2660, wire2661, wire2662, wire2663, wire2664, wire2665, wire2666, wire2667, wire2668, wire2669, wire2670, wire2671, wire2672, wire2673, wire2674, wire2675, wire2676, wire2677, wire2678, wire2679, wire2680, wire2681, wire2682, wire2683, wire2684, wire2685, wire2686, wire2687, wire2688, wire2689, wire2690, wire2691, wire2692, wire2693, wire2694, wire2695, wire2696, wire2697, wire2698, wire2699, wire2700, wire2701, wire2702, wire2703, wire2704, wire2705, wire2706, wire2707, wire2708, wire2709, wire2710, wire2711, wire2712, wire2713, wire2714, wire2715, wire2716, wire2717, wire2718, wire2719, wire2720, wire2721, wire2722, wire2723, wire2724, wire2725, wire2726, wire2727, wire2728, wire2729, wire2730, wire2731, wire2732, wire2733, wire2734, wire2735, wire2736, wire2737, wire2738, wire2739, wire2740, wire2741, wire2742, wire2743, wire2744, wire2745, wire2746, wire2747, wire2748, wire2749, wire2750, wire2751, wire2752, wire2753, wire2754, wire2755, wire2756, wire2757, wire2758, wire2759, wire2760, wire2761, wire2762, wire2763, wire2764, wire2765, wire2766, wire2767, wire2768, wire2769, wire2770, wire2771, wire2772, wire2773, wire2774, wire2775, wire2776, wire2777, wire2778, wire2779, wire2780, wire2781, wire2782, wire2783, wire2784, wire2785, wire2786, wire2787, wire2788, wire2789, wire2790, wire2791, wire2792, wire2793, wire2794, wire2795, wire2796, wire2797, wire2798, wire2799, wire2800, wire2801, wire2802, wire2803, wire2804, wire2805, wire2806, wire2807, wire2808, wire2809, wire2810, wire2811, wire2812, wire2813, wire2814, wire2815, wire2816, wire2817, wire2818, wire2819, wire2820, wire2821, wire2822, wire2823, wire2824, wire2825, wire2826, wire2827, wire2828, wire2829, wire2830, wire2831, wire2832, wire2833, wire2834, wire2835, wire2836, wire2837, wire2838, wire2839, wire2840, wire2841, wire2842, wire2843, wire2844, wire2845, wire2846, wire2847, wire2848, wire2849, wire2850, wire2851, wire2852, wire2853, wire2854, wire2855, wire2856, wire2857, wire2858, wire2859, wire2860, wire2861, wire2862, wire2863, wire2864, wire2865, wire2866, wire2867, wire2868, wire2869, wire2870, wire2871, wire2872, wire2873, wire2874, wire2875, wire2876, wire2877, wire2878, wire2879, wire2880, wire2881, wire2882, wire2883, wire2884, wire2885, wire2886, wire2887, wire2888, wire2889, wire2890, wire2891, wire2892, wire2893, wire2894, wire2895, wire2896, wire2897, wire2898, wire2899, wire2900, wire2901, wire2902, wire2903, wire2904, wire2905, wire2906, wire2907, wire2908, wire2909, wire2910, wire2911, wire2912, wire2913, wire2914, wire2915, wire2916, wire2917, wire2918, wire2919, wire2920, wire2921, wire2922, wire2923, wire2924, wire2925, wire2926, wire2927, wire2928, wire2929, wire2930, wire2931, wire2932, wire2933, wire2934, wire2935, wire2936, wire2937, wire2938, wire2939, wire2940, wire2941, wire2942, wire2943, wire2944, wire2945, wire2946, wire2947, wire2948, wire2949, wire2950, wire2951, wire2952, wire2953, wire2954, wire2955, wire2956, wire2957, wire2958, wire2959, wire2960, wire2961, wire2962, wire2963, wire2964, wire2965, wire2966, wire2967, wire2968, wire2969, wire2970, wire2971, wire2972, wire2973, wire2974, wire2975, wire2976, wire2977, wire2978, wire2979, wire2980, wire2981, wire2982, wire2983, wire2984, wire2985, wire2986, wire2987, wire2988, wire2989, wire2990, wire2991, wire2992, wire2993, wire2994, wire2995, wire2996, wire2997, wire2998, wire2999, wire3000, wire3001, wire3002, wire3003, wire3004, wire3005, wire3006, wire3007, wire3008, wire3009, wire3010, wire3011, wire3012, wire3013, wire3014, wire3015, wire3016, wire3017, wire3018, wire3019, wire3020, wire3021, wire3022, wire3023, wire3024, wire3025, wire3026, wire3027, wire3028, wire3029, wire3030, wire3031, wire3032, wire3033, wire3034, wire3035, wire3036, wire3037, wire3038, wire3039, wire3040, wire3041, wire3042, wire3043, wire3044, wire3045, wire3046, wire3047, wire3048, wire3049, wire3050, wire3051, wire3052, wire3053, wire3054, wire3055, wire3056, wire3057, wire3058, wire3059, wire3060, wire3061, wire3062, wire3063, wire3064, wire3065, wire3066, wire3067, wire3068, wire3069, wire3070, wire3071, wire3072, wire3073, wire3074, wire3075, wire3076, wire3077, wire3078, wire3079, wire3080, wire3081, wire3082, wire3083, wire3084, wire3085, wire3086, wire3087, wire3088, wire3089, wire3090, wire3091, wire3092, wire3093, wire3094, wire3095, wire3096, wire3097, wire3098, wire3099, wire3100, wire3101, wire3102, wire3103, wire3104, wire3105, wire3106, wire3107, wire3108, wire3109, wire3110, wire3111, wire3112, wire3113, wire3114, wire3115, wire3116, wire3117, wire3118, wire3119, wire3120, wire3121, wire3122, wire3123, wire3124, wire3125, wire3126, wire3127, wire3128, wire3129, wire3130, wire3131, wire3132, wire3133, wire3134, wire3135, wire3136, wire3137, wire3138, wire3139, wire3140, wire3141, wire3142, wire3143, wire3144, wire3145, wire3146, wire3147, wire3148, wire3149, wire3150, wire3151, wire3152, wire3153, wire3154, wire3155, wire3156, wire3157, wire3158, wire3159, wire3160, wire3161, wire3162, wire3163, wire3164, wire3165, wire3166, wire3167, wire3168, wire3169, wire3170, wire3171, wire3172, wire3173, wire3174, wire3175, wire3176, wire3177, wire3178, wire3179, wire3180, wire3181, wire3182, wire3183, wire3184, wire3185, wire3186, wire3187, wire3188, wire3189, wire3190, wire3191, wire3192, wire3193, wire3194, wire3195, wire3196, wire3197, wire3198, wire3199, wire3200, wire3201, wire3202, wire3203, wire3204, wire3205, wire3206, wire3207, wire3208, wire3209, wire3210, wire3211, wire3212, wire3213, wire3214, wire3215, wire3216, wire3217, wire3218, wire3219, wire3220, wire3221, wire3222, wire3223, wire3224, wire3225, wire3226, wire3227, wire3228, wire3229, wire3230, wire3231, wire3232, wire3233, wire3234, wire3235, wire3236, wire3237, wire3238, wire3239, wire3240, wire3241, wire3242, wire3243, wire3244, wire3245, wire3246, wire3247, wire3248, wire3249, wire3250, wire3251, wire3252, wire3253, wire3254, wire3255, wire3256, wire3257, wire3258, wire3259, wire3260, wire3261, wire3262, wire3263, wire3264, wire3265, wire3266, wire3267, wire3268, wire3269, wire3270, wire3271, wire3272, wire3273, wire3274, wire3275, wire3276, wire3277, wire3278, wire3279, wire3280, wire3281, wire3282, wire3283, wire3284, wire3285, wire3286, wire3287, wire3288, wire3289, wire3290, wire3291, wire3292, wire3293, wire3294, wire3295, wire3296, wire3297, wire3298, wire3299, wire3300, wire3301, wire3302, wire3303, wire3304, wire3305, wire3306, wire3307, wire3308, wire3309, wire3310, wire3311, wire3312, wire3313, wire3314, wire3315, wire3316, wire3317, wire3318, wire3319, wire3320, wire3321, wire3322, wire3323, wire3324, wire3325, wire3326, wire3327, wire3328, wire3329, wire3330, wire3331, wire3332, wire3333, wire3334, wire3335, wire3336, wire3337, wire3338, wire3339, wire3340, wire3341, wire3342, wire3343, wire3344, wire3345, wire3346, wire3347, wire3348, wire3349, wire3350, wire3351, wire3352, wire3353, wire3354, wire3355, wire3356, wire3357, wire3358, wire3359, wire3360, wire3361, wire3362, wire3363, wire3364, wire3365, wire3366, wire3367, wire3368, wire3369, wire3370, wire3371, wire3372, wire3373, wire3374, wire3375, wire3376, wire3377, wire3378, wire3379, wire3380, wire3381, wire3382, wire3383, wire3384, wire3385, wire3386, wire3387, wire3388, wire3389, wire3390, wire3391, wire3392, wire3393, wire3394, wire3395, wire3396, wire3397, wire3398, wire3399, wire3400, wire3401, wire3402, wire3403, wire3404, wire3405, wire3406, wire3407, wire3408, wire3409, wire3410, wire3411, wire3412, wire3413, wire3414, wire3415, wire3416, wire3417, wire3418, wire3419, wire3420, wire3421, wire3422, wire3423, wire3424, wire3425, wire3426, wire3427, wire3428, wire3429, wire3430, wire3431, wire3432, wire3433, wire3434, wire3435, wire3436, wire3437, wire3438, wire3439, wire3440, wire3441, wire3442, wire3443, wire3444, wire3445, wire3446, wire3447, wire3448, wire3449, wire3450, wire3451, wire3452, wire3453, wire3454, wire3455, wire3456, wire3457, wire3458, wire3459, wire3460, wire3461, wire3462, wire3463, wire3464, wire3465, wire3466, wire3467, wire3468, wire3469, wire3470, wire3471, wire3472, wire3473, wire3474, wire3475, wire3476, wire3477, wire3478, wire3479, wire3480, wire3481, wire3482, wire3483, wire3484, wire3485, wire3486, wire3487, wire3488, wire3489, wire3490, wire3491, wire3492, wire3493, wire3494, wire3495, wire3496, wire3497, wire3498, wire3499, wire3500, wire3501, wire3502, wire3503, wire3504, wire3505, wire3506, wire3507, wire3508, wire3509, wire3510, wire3511, wire3512, wire3513, wire3514, wire3515, wire3516, wire3517, wire3518, wire3519, wire3520, wire3521, wire3522, wire3523, wire3524, wire3525, wire3526, wire3527, wire3528, wire3529, wire3530, wire3531, wire3532, wire3533, wire3534, wire3535, wire3536, wire3537, wire3538, wire3539, wire3540, wire3541, wire3542, wire3543, wire3544, wire3545, wire3546, wire3547, wire3548, wire3549, wire3550, wire3551, wire3552, wire3553, wire3554, wire3555, wire3556, wire3557, wire3558, wire3559, wire3560, wire3561, wire3562, wire3563, wire3564, wire3565, wire3566, wire3567, wire3568, wire3569, wire3570, wire3571, wire3572, wire3573, wire3574, wire3575, wire3576, wire3577, wire3578, wire3579, wire3580, wire3581, wire3582, wire3583, wire3584, wire3585, wire3586, wire3587, wire3588, wire3589, wire3590, wire3591, wire3592, wire3593, wire3594, wire3595, wire3596, wire3597, wire3598, wire3599, wire3600, wire3601, wire3602, wire3603, wire3604, wire3605, wire3606, wire3607, wire3608, wire3609, wire3610, wire3611, wire3612, wire3613, wire3614, wire3615, wire3616, wire3617, wire3618, wire3619, wire3620, wire3621, wire3622, wire3623, wire3624, wire3625, wire3626, wire3627, wire3628, wire3629, wire3630, wire3631, wire3632, wire3633, wire3634, wire3635, wire3636, wire3637, wire3638, wire3639, wire3640, wire3641, wire3642, wire3643, wire3644, wire3645, wire3646, wire3647, wire3648, wire3649, wire3650, wire3651, wire3652, wire3653, wire3654, wire3655, wire3656, wire3657, wire3658, wire3659, wire3660, wire3661, wire3662, wire3663, wire3664, wire3665, wire3666, wire3667, wire3668, wire3669, wire3670, wire3671, wire3672, wire3673, wire3674, wire3675, wire3676, wire3677, wire3678, wire3679, wire3680, wire3681, wire3682, wire3683, wire3684, wire3685, wire3686, wire3687, wire3688, wire3689, wire3690, wire3691, wire3692, wire3693, wire3694, wire3695, wire3696, wire3697, wire3698, wire3699, wire3700, wire3701, wire3702, wire3703, wire3704, wire3705, wire3706, wire3707, wire3708, wire3709, wire3710, wire3711, wire3712, wire3713, wire3714, wire3715, wire3716, wire3717, wire3718, wire3719, wire3720, wire3721, wire3722, wire3723, wire3724, wire3725, wire3726, wire3727, wire3728, wire3729, wire3730, wire3731, wire3732, wire3733, wire3734, wire3735, wire3736, wire3737, wire3738, wire3739, wire3740, wire3741, wire3742, wire3743, wire3744, wire3745, wire3746, wire3747, wire3748, wire3749, wire3750, wire3751, wire3752, wire3753, wire3754, wire3755, wire3756, wire3757, wire3758, wire3759, wire3760, wire3761, wire3762, wire3763, wire3764, wire3765, wire3766, wire3767, wire3768, wire3769, wire3770, wire3771, wire3772, wire3773, wire3774, wire3775, wire3776, wire3777, wire3778, wire3779, wire3780, wire3781, wire3782, wire3783, wire3784, wire3785, wire3786, wire3787, wire3788, wire3789, wire3790, wire3791, wire3792, wire3793, wire3794, wire3795, wire3796, wire3797, wire3798, wire3799, wire3800, wire3801, wire3802, wire3803, wire3804, wire3805, wire3806, wire3807, wire3808, wire3809, wire3810, wire3811, wire3812, wire3813, wire3814, wire3815, wire3816, wire3817, wire3818, wire3819, wire3820, wire3821, wire3822, wire3823, wire3824, wire3825, wire3826, wire3827, wire3828, wire3829, wire3830, wire3831, wire3832, wire3833, wire3834, wire3835, wire3836, wire3837, wire3838, wire3839, wire3840, wire3841, wire3842, wire3843, wire3844, wire3845, wire3846, wire3847, wire3848, wire3849, wire3850, wire3851, wire3852, wire3853, wire3854, wire3855, wire3856, wire3857, wire3858, wire3859, wire3860, wire3861, wire3862, wire3863, wire3864, wire3865, wire3866, wire3867, wire3868, wire3869, wire3870, wire3871, wire3872, wire3873, wire3874, wire3875, wire3876, wire3877, wire3878, wire3879, wire3880, wire3881, wire3882, wire3883, wire3884, wire3885, wire3886, wire3887, wire3888, wire3889, wire3890, wire3891, wire3892, wire3893, wire3894, wire3895, wire3896, wire3897, wire3898, wire3899, wire3900, wire3901, wire3902, wire3903, wire3904, wire3905, wire3906, wire3907, wire3908, wire3909, wire3910, wire3911, wire3912, wire3913, wire3914, wire3915, wire3916, wire3917, wire3918, wire3919, wire3920, wire3921, wire3922, wire3923, wire3924, wire3925, wire3926, wire3927, wire3928, wire3929, wire3930, wire3931, wire3932, wire3933, wire3934, wire3935, wire3936, wire3937, wire3938, wire3939, wire3940, wire3941, wire3942, wire3943, wire3944, wire3945, wire3946, wire3947, wire3948, wire3949, wire3950, wire3951, wire3952, wire3953, wire3954, wire3955, wire3956, wire3957, wire3958, wire3959, wire3960, wire3961, wire3962, wire3963, wire3964, wire3965, wire3966, wire3967, wire3968, wire3969, wire3970, wire3971, wire3972, wire3973, wire3974, wire3975, wire3976, wire3977, wire3978, wire3979, wire3980, wire3981, wire3982, wire3983, wire3984, wire3985, wire3986, wire3987, wire3988, wire3989, wire3990, wire3991, wire3992, wire3993, wire3994, wire3995, wire3996, wire3997, wire3998, wire3999, wire4000, wire4001, wire4002, wire4003, wire4004, wire4005, wire4006, wire4007, wire4008, wire4009, wire4010, wire4011, wire4012, wire4013, wire4014, wire4015, wire4016, wire4017, wire4018, wire4019, wire4020, wire4021, wire4022, wire4023, wire4024, wire4025, wire4026, wire4027, wire4028, wire4029, wire4030, wire4031, wire4032, wire4033, wire4034, wire4035, wire4036, wire4037, wire4038, wire4039, wire4040, wire4041, wire4042, wire4043, wire4044, wire4045, wire4046, wire4047, wire4048, wire4049, wire4050, wire4051, wire4052, wire4053, wire4054, wire4055, wire4056, wire4057, wire4058, wire4059, wire4060, wire4061, wire4062, wire4063, wire4064, wire4065, wire4066, wire4067, wire4068, wire4069, wire4070, wire4071, wire4072, wire4073, wire4074, wire4075, wire4076, wire4077, wire4078, wire4079, wire4080, wire4081, wire4082, wire4083, wire4084, wire4085, wire4086, wire4087, wire4088, wire4089, wire4090, wire4091, wire4092, wire4093, wire4094, wire4095;
    assign wire0 = {5'd2, 5'd1};
    assign wire1 = {5'd2, 5'd1};
    assign wire2 = {5'd2, 5'd1};
    assign wire3 = {5'd2, 5'd1};
    assign wire4 = {5'd2, 5'd1};
    assign wire5 = {5'd2, 5'd1};
    assign wire6 = {5'd2, 5'd1};
    assign wire7 = {5'd2, 5'd1};
    assign wire8 = {5'd2, 5'd1};
    assign wire9 = {5'd2, 5'd1};
    assign wire10 = {5'd2, 5'd1};
    assign wire11 = {5'd2, 5'd1};
    assign wire12 = {5'd2, 5'd1};
    assign wire13 = {5'd2, 5'd1};
    assign wire14 = {5'd2, 5'd1};
    assign wire15 = {5'd2, 5'd1};
    assign wire16 = {5'd2, 5'd1};
    assign wire17 = {5'd2, 5'd1};
    assign wire18 = {5'd2, 5'd1};
    assign wire19 = {5'd2, 5'd1};
    assign wire20 = {5'd2, 5'd1};
    assign wire21 = {5'd2, 5'd1};
    assign wire22 = {5'd2, 5'd1};
    assign wire23 = {5'd2, 5'd1};
    assign wire24 = {5'd2, 5'd1};
    assign wire25 = {5'd2, 5'd1};
    assign wire26 = {5'd2, 5'd1};
    assign wire27 = {5'd2, 5'd1};
    assign wire28 = {5'd2, 5'd1};
    assign wire29 = {5'd2, 5'd1};
    assign wire30 = {5'd2, 5'd1};
    assign wire31 = {5'd2, 5'd1};
    assign wire32 = {5'd3, 5'd1};
    assign wire33 = {5'd3, 5'd1};
    assign wire34 = {5'd3, 5'd1};
    assign wire35 = {5'd3, 5'd1};
    assign wire36 = {5'd3, 5'd1};
    assign wire37 = {5'd3, 5'd1};
    assign wire38 = {5'd3, 5'd1};
    assign wire39 = {5'd3, 5'd1};
    assign wire40 = {5'd3, 5'd1};
    assign wire41 = {5'd3, 5'd1};
    assign wire42 = {5'd3, 5'd1};
    assign wire43 = {5'd3, 5'd1};
    assign wire44 = {5'd3, 5'd1};
    assign wire45 = {5'd3, 5'd1};
    assign wire46 = {5'd3, 5'd1};
    assign wire47 = {5'd3, 5'd1};
    assign wire48 = {5'd3, 5'd1};
    assign wire49 = {5'd3, 5'd1};
    assign wire50 = {5'd3, 5'd1};
    assign wire51 = {5'd3, 5'd1};
    assign wire52 = {5'd3, 5'd1};
    assign wire53 = {5'd3, 5'd1};
    assign wire54 = {5'd3, 5'd1};
    assign wire55 = {5'd3, 5'd1};
    assign wire56 = {5'd3, 5'd1};
    assign wire57 = {5'd3, 5'd1};
    assign wire58 = {5'd3, 5'd1};
    assign wire59 = {5'd3, 5'd1};
    assign wire60 = {5'd3, 5'd1};
    assign wire61 = {5'd3, 5'd1};
    assign wire62 = {5'd3, 5'd1};
    assign wire63 = {5'd3, 5'd1};
    assign wire64 = {5'd5, 5'd1};
    assign wire65 = {5'd5, 5'd1};
    assign wire66 = {5'd5, 5'd1};
    assign wire67 = {5'd5, 5'd1};
    assign wire68 = {5'd5, 5'd1};
    assign wire69 = {5'd5, 5'd1};
    assign wire70 = {5'd5, 5'd1};
    assign wire71 = {5'd5, 5'd1};
    assign wire72 = {5'd5, 5'd1};
    assign wire73 = {5'd5, 5'd1};
    assign wire74 = {5'd5, 5'd1};
    assign wire75 = {5'd5, 5'd1};
    assign wire76 = {5'd5, 5'd1};
    assign wire77 = {5'd5, 5'd1};
    assign wire78 = {5'd5, 5'd1};
    assign wire79 = {5'd5, 5'd1};
    assign wire80 = {5'd5, 5'd1};
    assign wire81 = {5'd5, 5'd1};
    assign wire82 = {5'd5, 5'd1};
    assign wire83 = {5'd5, 5'd1};
    assign wire84 = {5'd5, 5'd1};
    assign wire85 = {5'd5, 5'd1};
    assign wire86 = {5'd5, 5'd1};
    assign wire87 = {5'd5, 5'd1};
    assign wire88 = {5'd5, 5'd1};
    assign wire89 = {5'd5, 5'd1};
    assign wire90 = {5'd5, 5'd1};
    assign wire91 = {5'd5, 5'd1};
    assign wire92 = {5'd5, 5'd1};
    assign wire93 = {5'd5, 5'd1};
    assign wire94 = {5'd5, 5'd1};
    assign wire95 = {5'd5, 5'd1};
    assign wire96 = {5'd7, 5'd1};
    assign wire97 = {5'd7, 5'd1};
    assign wire98 = {5'd7, 5'd1};
    assign wire99 = {5'd7, 5'd1};
    assign wire100 = {5'd7, 5'd1};
    assign wire101 = {5'd7, 5'd1};
    assign wire102 = {5'd7, 5'd1};
    assign wire103 = {5'd7, 5'd1};
    assign wire104 = {5'd7, 5'd1};
    assign wire105 = {5'd7, 5'd1};
    assign wire106 = {5'd7, 5'd1};
    assign wire107 = {5'd7, 5'd1};
    assign wire108 = {5'd7, 5'd1};
    assign wire109 = {5'd7, 5'd1};
    assign wire110 = {5'd7, 5'd1};
    assign wire111 = {5'd7, 5'd1};
    assign wire112 = {5'd7, 5'd1};
    assign wire113 = {5'd7, 5'd1};
    assign wire114 = {5'd7, 5'd1};
    assign wire115 = {5'd7, 5'd1};
    assign wire116 = {5'd7, 5'd1};
    assign wire117 = {5'd7, 5'd1};
    assign wire118 = {5'd7, 5'd1};
    assign wire119 = {5'd7, 5'd1};
    assign wire120 = {5'd7, 5'd1};
    assign wire121 = {5'd7, 5'd1};
    assign wire122 = {5'd7, 5'd1};
    assign wire123 = {5'd7, 5'd1};
    assign wire124 = {5'd7, 5'd1};
    assign wire125 = {5'd7, 5'd1};
    assign wire126 = {5'd7, 5'd1};
    assign wire127 = {5'd7, 5'd1};
    assign wire128 = {5'd3, 5'd2};
    assign wire129 = {5'd3, 5'd2};
    assign wire130 = {5'd3, 5'd2};
    assign wire131 = {5'd3, 5'd2};
    assign wire132 = {5'd4, 5'd3};
    assign wire133 = {5'd7, 5'd6};
    assign wire134 = {5'd3, 5'd2};
    assign wire135 = {5'd3, 5'd2};
    assign wire136 = {5'd4, 5'd3};
    assign wire137 = {5'd4, 5'd3};
    assign wire138 = {5'd4, 5'd3};
    assign wire139 = {5'd4, 5'd3};
    assign wire140 = {5'd5, 5'd4};
    assign wire141 = {5'd4, 5'd3};
    assign wire142 = {5'd4, 5'd3};
    assign wire143 = {5'd4, 5'd3};
    assign wire144 = {5'd7, 5'd6};
    assign wire145 = {5'd7, 5'd6};
    assign wire146 = {5'd7, 5'd6};
    assign wire147 = {5'd7, 5'd6};
    assign wire148 = {5'd8, 5'd7};
    assign wire149 = {5'd7, 5'd6};
    assign wire150 = {5'd7, 5'd6};
    assign wire151 = {5'd7, 5'd6};
    assign wire152 = {5'd3, 5'd2};
    assign wire153 = {5'd3, 5'd2};
    assign wire154 = {5'd3, 5'd2};
    assign wire155 = {5'd3, 5'd2};
    assign wire156 = {5'd3, 5'd2};
    assign wire157 = {5'd3, 5'd2};
    assign wire158 = {5'd3, 5'd2};
    assign wire159 = {5'd3, 5'd2};
    assign wire160 = {5'd4, 5'd2};
    assign wire161 = {5'd4, 5'd2};
    assign wire162 = {5'd4, 5'd2};
    assign wire163 = {5'd4, 5'd2};
    assign wire164 = {5'd5, 5'd3};
    assign wire165 = {5'd8, 5'd6};
    assign wire166 = {5'd4, 5'd2};
    assign wire167 = {5'd4, 5'd2};
    assign wire168 = {5'd5, 5'd3};
    assign wire169 = {5'd5, 5'd3};
    assign wire170 = {5'd5, 5'd3};
    assign wire171 = {5'd5, 5'd3};
    assign wire172 = {5'd6, 5'd4};
    assign wire173 = {5'd5, 5'd3};
    assign wire174 = {5'd5, 5'd3};
    assign wire175 = {5'd5, 5'd3};
    assign wire176 = {5'd8, 5'd6};
    assign wire177 = {5'd8, 5'd6};
    assign wire178 = {5'd8, 5'd6};
    assign wire179 = {5'd8, 5'd6};
    assign wire180 = {5'd9, 5'd7};
    assign wire181 = {5'd8, 5'd6};
    assign wire182 = {5'd8, 5'd6};
    assign wire183 = {5'd8, 5'd6};
    assign wire184 = {5'd4, 5'd2};
    assign wire185 = {5'd4, 5'd2};
    assign wire186 = {5'd4, 5'd2};
    assign wire187 = {5'd4, 5'd2};
    assign wire188 = {5'd4, 5'd2};
    assign wire189 = {5'd4, 5'd2};
    assign wire190 = {5'd4, 5'd2};
    assign wire191 = {5'd4, 5'd2};
    assign wire192 = {5'd6, 5'd2};
    assign wire193 = {5'd6, 5'd2};
    assign wire194 = {5'd6, 5'd2};
    assign wire195 = {5'd6, 5'd2};
    assign wire196 = {5'd7, 5'd3};
    assign wire197 = {5'd10, 5'd6};
    assign wire198 = {5'd6, 5'd2};
    assign wire199 = {5'd6, 5'd2};
    assign wire200 = {5'd7, 5'd3};
    assign wire201 = {5'd7, 5'd3};
    assign wire202 = {5'd7, 5'd3};
    assign wire203 = {5'd7, 5'd3};
    assign wire204 = {5'd8, 5'd4};
    assign wire205 = {5'd7, 5'd3};
    assign wire206 = {5'd7, 5'd3};
    assign wire207 = {5'd7, 5'd3};
    assign wire208 = {5'd10, 5'd6};
    assign wire209 = {5'd10, 5'd6};
    assign wire210 = {5'd10, 5'd6};
    assign wire211 = {5'd10, 5'd6};
    assign wire212 = {5'd11, 5'd7};
    assign wire213 = {5'd10, 5'd6};
    assign wire214 = {5'd10, 5'd6};
    assign wire215 = {5'd10, 5'd6};
    assign wire216 = {5'd6, 5'd2};
    assign wire217 = {5'd6, 5'd2};
    assign wire218 = {5'd6, 5'd2};
    assign wire219 = {5'd6, 5'd2};
    assign wire220 = {5'd6, 5'd2};
    assign wire221 = {5'd6, 5'd2};
    assign wire222 = {5'd6, 5'd2};
    assign wire223 = {5'd6, 5'd2};
    assign wire224 = {5'd8, 5'd2};
    assign wire225 = {5'd8, 5'd2};
    assign wire226 = {5'd8, 5'd2};
    assign wire227 = {5'd8, 5'd2};
    assign wire228 = {5'd9, 5'd3};
    assign wire229 = {5'd12, 5'd6};
    assign wire230 = {5'd8, 5'd2};
    assign wire231 = {5'd8, 5'd2};
    assign wire232 = {5'd9, 5'd3};
    assign wire233 = {5'd9, 5'd3};
    assign wire234 = {5'd9, 5'd3};
    assign wire235 = {5'd9, 5'd3};
    assign wire236 = {5'd10, 5'd4};
    assign wire237 = {5'd9, 5'd3};
    assign wire238 = {5'd9, 5'd3};
    assign wire239 = {5'd9, 5'd3};
    assign wire240 = {5'd12, 5'd6};
    assign wire241 = {5'd12, 5'd6};
    assign wire242 = {5'd12, 5'd6};
    assign wire243 = {5'd12, 5'd6};
    assign wire244 = {5'd13, 5'd7};
    assign wire245 = {5'd12, 5'd6};
    assign wire246 = {5'd12, 5'd6};
    assign wire247 = {5'd12, 5'd6};
    assign wire248 = {5'd8, 5'd2};
    assign wire249 = {5'd8, 5'd2};
    assign wire250 = {5'd8, 5'd2};
    assign wire251 = {5'd8, 5'd2};
    assign wire252 = {5'd8, 5'd2};
    assign wire253 = {5'd8, 5'd2};
    assign wire254 = {5'd8, 5'd2};
    assign wire255 = {5'd8, 5'd2};
    assign wire256 = {5'd3, 5'd2};
    assign wire257 = {5'd3, 5'd2};
    assign wire258 = {5'd3, 5'd2};
    assign wire259 = {5'd3, 5'd2};
    assign wire260 = {5'd3, 5'd2};
    assign wire261 = {5'd3, 5'd2};
    assign wire262 = {5'd3, 5'd2};
    assign wire263 = {5'd3, 5'd2};
    assign wire264 = {5'd3, 5'd2};
    assign wire265 = {5'd3, 5'd2};
    assign wire266 = {5'd3, 5'd2};
    assign wire267 = {5'd3, 5'd2};
    assign wire268 = {5'd3, 5'd2};
    assign wire269 = {5'd3, 5'd2};
    assign wire270 = {5'd3, 5'd2};
    assign wire271 = {5'd3, 5'd2};
    assign wire272 = {5'd3, 5'd2};
    assign wire273 = {5'd3, 5'd2};
    assign wire274 = {5'd3, 5'd2};
    assign wire275 = {5'd3, 5'd2};
    assign wire276 = {5'd3, 5'd2};
    assign wire277 = {5'd3, 5'd2};
    assign wire278 = {5'd3, 5'd2};
    assign wire279 = {5'd3, 5'd2};
    assign wire280 = {5'd3, 5'd2};
    assign wire281 = {5'd3, 5'd2};
    assign wire282 = {5'd3, 5'd2};
    assign wire283 = {5'd3, 5'd2};
    assign wire284 = {5'd3, 5'd2};
    assign wire285 = {5'd3, 5'd2};
    assign wire286 = {5'd3, 5'd2};
    assign wire287 = {5'd3, 5'd2};
    assign wire288 = {5'd4, 5'd2};
    assign wire289 = {5'd4, 5'd2};
    assign wire290 = {5'd4, 5'd2};
    assign wire291 = {5'd4, 5'd2};
    assign wire292 = {5'd4, 5'd2};
    assign wire293 = {5'd4, 5'd2};
    assign wire294 = {5'd4, 5'd2};
    assign wire295 = {5'd4, 5'd2};
    assign wire296 = {5'd4, 5'd2};
    assign wire297 = {5'd4, 5'd2};
    assign wire298 = {5'd4, 5'd2};
    assign wire299 = {5'd4, 5'd2};
    assign wire300 = {5'd4, 5'd2};
    assign wire301 = {5'd4, 5'd2};
    assign wire302 = {5'd4, 5'd2};
    assign wire303 = {5'd4, 5'd2};
    assign wire304 = {5'd4, 5'd2};
    assign wire305 = {5'd4, 5'd2};
    assign wire306 = {5'd4, 5'd2};
    assign wire307 = {5'd4, 5'd2};
    assign wire308 = {5'd4, 5'd2};
    assign wire309 = {5'd4, 5'd2};
    assign wire310 = {5'd4, 5'd2};
    assign wire311 = {5'd4, 5'd2};
    assign wire312 = {5'd4, 5'd2};
    assign wire313 = {5'd4, 5'd2};
    assign wire314 = {5'd4, 5'd2};
    assign wire315 = {5'd4, 5'd2};
    assign wire316 = {5'd4, 5'd2};
    assign wire317 = {5'd4, 5'd2};
    assign wire318 = {5'd4, 5'd2};
    assign wire319 = {5'd4, 5'd2};
    assign wire320 = {5'd6, 5'd2};
    assign wire321 = {5'd6, 5'd2};
    assign wire322 = {5'd6, 5'd2};
    assign wire323 = {5'd6, 5'd2};
    assign wire324 = {5'd6, 5'd2};
    assign wire325 = {5'd6, 5'd2};
    assign wire326 = {5'd6, 5'd2};
    assign wire327 = {5'd6, 5'd2};
    assign wire328 = {5'd6, 5'd2};
    assign wire329 = {5'd6, 5'd2};
    assign wire330 = {5'd6, 5'd2};
    assign wire331 = {5'd6, 5'd2};
    assign wire332 = {5'd6, 5'd2};
    assign wire333 = {5'd6, 5'd2};
    assign wire334 = {5'd6, 5'd2};
    assign wire335 = {5'd6, 5'd2};
    assign wire336 = {5'd6, 5'd2};
    assign wire337 = {5'd6, 5'd2};
    assign wire338 = {5'd6, 5'd2};
    assign wire339 = {5'd6, 5'd2};
    assign wire340 = {5'd6, 5'd2};
    assign wire341 = {5'd6, 5'd2};
    assign wire342 = {5'd6, 5'd2};
    assign wire343 = {5'd6, 5'd2};
    assign wire344 = {5'd6, 5'd2};
    assign wire345 = {5'd6, 5'd2};
    assign wire346 = {5'd6, 5'd2};
    assign wire347 = {5'd6, 5'd2};
    assign wire348 = {5'd6, 5'd2};
    assign wire349 = {5'd6, 5'd2};
    assign wire350 = {5'd6, 5'd2};
    assign wire351 = {5'd6, 5'd2};
    assign wire352 = {5'd8, 5'd2};
    assign wire353 = {5'd8, 5'd2};
    assign wire354 = {5'd8, 5'd2};
    assign wire355 = {5'd8, 5'd2};
    assign wire356 = {5'd8, 5'd2};
    assign wire357 = {5'd8, 5'd2};
    assign wire358 = {5'd8, 5'd2};
    assign wire359 = {5'd8, 5'd2};
    assign wire360 = {5'd8, 5'd2};
    assign wire361 = {5'd8, 5'd2};
    assign wire362 = {5'd8, 5'd2};
    assign wire363 = {5'd8, 5'd2};
    assign wire364 = {5'd8, 5'd2};
    assign wire365 = {5'd8, 5'd2};
    assign wire366 = {5'd8, 5'd2};
    assign wire367 = {5'd8, 5'd2};
    assign wire368 = {5'd8, 5'd2};
    assign wire369 = {5'd8, 5'd2};
    assign wire370 = {5'd8, 5'd2};
    assign wire371 = {5'd8, 5'd2};
    assign wire372 = {5'd8, 5'd2};
    assign wire373 = {5'd8, 5'd2};
    assign wire374 = {5'd8, 5'd2};
    assign wire375 = {5'd8, 5'd2};
    assign wire376 = {5'd8, 5'd2};
    assign wire377 = {5'd8, 5'd2};
    assign wire378 = {5'd8, 5'd2};
    assign wire379 = {5'd8, 5'd2};
    assign wire380 = {5'd8, 5'd2};
    assign wire381 = {5'd8, 5'd2};
    assign wire382 = {5'd8, 5'd2};
    assign wire383 = {5'd8, 5'd2};
    assign wire384 = {5'd4, 5'd3};
    assign wire385 = {5'd4, 5'd3};
    assign wire386 = {5'd4, 5'd3};
    assign wire387 = {5'd4, 5'd3};
    assign wire388 = {5'd5, 5'd4};
    assign wire389 = {5'd8, 5'd7};
    assign wire390 = {5'd4, 5'd3};
    assign wire391 = {5'd4, 5'd3};
    assign wire392 = {5'd5, 5'd4};
    assign wire393 = {5'd5, 5'd4};
    assign wire394 = {5'd5, 5'd4};
    assign wire395 = {5'd5, 5'd4};
    assign wire396 = {5'd6, 5'd5};
    assign wire397 = {5'd5, 5'd4};
    assign wire398 = {5'd5, 5'd4};
    assign wire399 = {5'd5, 5'd4};
    assign wire400 = {5'd8, 5'd7};
    assign wire401 = {5'd8, 5'd7};
    assign wire402 = {5'd8, 5'd7};
    assign wire403 = {5'd8, 5'd7};
    assign wire404 = {5'd9, 5'd8};
    assign wire405 = {5'd8, 5'd7};
    assign wire406 = {5'd8, 5'd7};
    assign wire407 = {5'd8, 5'd7};
    assign wire408 = {5'd4, 5'd3};
    assign wire409 = {5'd4, 5'd3};
    assign wire410 = {5'd4, 5'd3};
    assign wire411 = {5'd4, 5'd3};
    assign wire412 = {5'd4, 5'd3};
    assign wire413 = {5'd4, 5'd3};
    assign wire414 = {5'd4, 5'd3};
    assign wire415 = {5'd4, 5'd3};
    assign wire416 = {5'd5, 5'd3};
    assign wire417 = {5'd5, 5'd3};
    assign wire418 = {5'd5, 5'd3};
    assign wire419 = {5'd5, 5'd3};
    assign wire420 = {5'd6, 5'd4};
    assign wire421 = {5'd9, 5'd7};
    assign wire422 = {5'd5, 5'd3};
    assign wire423 = {5'd5, 5'd3};
    assign wire424 = {5'd6, 5'd4};
    assign wire425 = {5'd6, 5'd4};
    assign wire426 = {5'd6, 5'd4};
    assign wire427 = {5'd6, 5'd4};
    assign wire428 = {5'd7, 5'd5};
    assign wire429 = {5'd6, 5'd4};
    assign wire430 = {5'd6, 5'd4};
    assign wire431 = {5'd6, 5'd4};
    assign wire432 = {5'd9, 5'd7};
    assign wire433 = {5'd9, 5'd7};
    assign wire434 = {5'd9, 5'd7};
    assign wire435 = {5'd9, 5'd7};
    assign wire436 = {5'd10, 5'd8};
    assign wire437 = {5'd9, 5'd7};
    assign wire438 = {5'd9, 5'd7};
    assign wire439 = {5'd9, 5'd7};
    assign wire440 = {5'd5, 5'd3};
    assign wire441 = {5'd5, 5'd3};
    assign wire442 = {5'd5, 5'd3};
    assign wire443 = {5'd5, 5'd3};
    assign wire444 = {5'd5, 5'd3};
    assign wire445 = {5'd5, 5'd3};
    assign wire446 = {5'd5, 5'd3};
    assign wire447 = {5'd5, 5'd3};
    assign wire448 = {5'd7, 5'd3};
    assign wire449 = {5'd7, 5'd3};
    assign wire450 = {5'd7, 5'd3};
    assign wire451 = {5'd7, 5'd3};
    assign wire452 = {5'd8, 5'd4};
    assign wire453 = {5'd11, 5'd7};
    assign wire454 = {5'd7, 5'd3};
    assign wire455 = {5'd7, 5'd3};
    assign wire456 = {5'd8, 5'd4};
    assign wire457 = {5'd8, 5'd4};
    assign wire458 = {5'd8, 5'd4};
    assign wire459 = {5'd8, 5'd4};
    assign wire460 = {5'd9, 5'd5};
    assign wire461 = {5'd8, 5'd4};
    assign wire462 = {5'd8, 5'd4};
    assign wire463 = {5'd8, 5'd4};
    assign wire464 = {5'd11, 5'd7};
    assign wire465 = {5'd11, 5'd7};
    assign wire466 = {5'd11, 5'd7};
    assign wire467 = {5'd11, 5'd7};
    assign wire468 = {5'd12, 5'd8};
    assign wire469 = {5'd11, 5'd7};
    assign wire470 = {5'd11, 5'd7};
    assign wire471 = {5'd11, 5'd7};
    assign wire472 = {5'd7, 5'd3};
    assign wire473 = {5'd7, 5'd3};
    assign wire474 = {5'd7, 5'd3};
    assign wire475 = {5'd7, 5'd3};
    assign wire476 = {5'd7, 5'd3};
    assign wire477 = {5'd7, 5'd3};
    assign wire478 = {5'd7, 5'd3};
    assign wire479 = {5'd7, 5'd3};
    assign wire480 = {5'd9, 5'd3};
    assign wire481 = {5'd9, 5'd3};
    assign wire482 = {5'd9, 5'd3};
    assign wire483 = {5'd9, 5'd3};
    assign wire484 = {5'd10, 5'd4};
    assign wire485 = {5'd13, 5'd7};
    assign wire486 = {5'd9, 5'd3};
    assign wire487 = {5'd9, 5'd3};
    assign wire488 = {5'd10, 5'd4};
    assign wire489 = {5'd10, 5'd4};
    assign wire490 = {5'd10, 5'd4};
    assign wire491 = {5'd10, 5'd4};
    assign wire492 = {5'd11, 5'd5};
    assign wire493 = {5'd10, 5'd4};
    assign wire494 = {5'd10, 5'd4};
    assign wire495 = {5'd10, 5'd4};
    assign wire496 = {5'd13, 5'd7};
    assign wire497 = {5'd13, 5'd7};
    assign wire498 = {5'd13, 5'd7};
    assign wire499 = {5'd13, 5'd7};
    assign wire500 = {5'd14, 5'd8};
    assign wire501 = {5'd13, 5'd7};
    assign wire502 = {5'd13, 5'd7};
    assign wire503 = {5'd13, 5'd7};
    assign wire504 = {5'd9, 5'd3};
    assign wire505 = {5'd9, 5'd3};
    assign wire506 = {5'd9, 5'd3};
    assign wire507 = {5'd9, 5'd3};
    assign wire508 = {5'd9, 5'd3};
    assign wire509 = {5'd9, 5'd3};
    assign wire510 = {5'd9, 5'd3};
    assign wire511 = {5'd9, 5'd3};
    assign wire512 = {5'd3, 5'd2};
    assign wire513 = {5'd3, 5'd2};
    assign wire514 = {5'd3, 5'd2};
    assign wire515 = {5'd3, 5'd2};
    assign wire516 = {5'd3, 5'd2};
    assign wire517 = {5'd3, 5'd2};
    assign wire518 = {5'd3, 5'd2};
    assign wire519 = {5'd3, 5'd2};
    assign wire520 = {5'd3, 5'd2};
    assign wire521 = {5'd3, 5'd2};
    assign wire522 = {5'd3, 5'd2};
    assign wire523 = {5'd3, 5'd2};
    assign wire524 = {5'd3, 5'd2};
    assign wire525 = {5'd3, 5'd2};
    assign wire526 = {5'd3, 5'd2};
    assign wire527 = {5'd3, 5'd2};
    assign wire528 = {5'd3, 5'd2};
    assign wire529 = {5'd3, 5'd2};
    assign wire530 = {5'd3, 5'd2};
    assign wire531 = {5'd3, 5'd2};
    assign wire532 = {5'd3, 5'd2};
    assign wire533 = {5'd3, 5'd2};
    assign wire534 = {5'd3, 5'd2};
    assign wire535 = {5'd3, 5'd2};
    assign wire536 = {5'd3, 5'd2};
    assign wire537 = {5'd3, 5'd2};
    assign wire538 = {5'd3, 5'd2};
    assign wire539 = {5'd3, 5'd2};
    assign wire540 = {5'd3, 5'd2};
    assign wire541 = {5'd3, 5'd2};
    assign wire542 = {5'd3, 5'd2};
    assign wire543 = {5'd3, 5'd2};
    assign wire544 = {5'd4, 5'd2};
    assign wire545 = {5'd4, 5'd2};
    assign wire546 = {5'd4, 5'd2};
    assign wire547 = {5'd4, 5'd2};
    assign wire548 = {5'd4, 5'd2};
    assign wire549 = {5'd4, 5'd2};
    assign wire550 = {5'd4, 5'd2};
    assign wire551 = {5'd4, 5'd2};
    assign wire552 = {5'd4, 5'd2};
    assign wire553 = {5'd4, 5'd2};
    assign wire554 = {5'd4, 5'd2};
    assign wire555 = {5'd4, 5'd2};
    assign wire556 = {5'd4, 5'd2};
    assign wire557 = {5'd4, 5'd2};
    assign wire558 = {5'd4, 5'd2};
    assign wire559 = {5'd4, 5'd2};
    assign wire560 = {5'd4, 5'd2};
    assign wire561 = {5'd4, 5'd2};
    assign wire562 = {5'd4, 5'd2};
    assign wire563 = {5'd4, 5'd2};
    assign wire564 = {5'd4, 5'd2};
    assign wire565 = {5'd4, 5'd2};
    assign wire566 = {5'd4, 5'd2};
    assign wire567 = {5'd4, 5'd2};
    assign wire568 = {5'd4, 5'd2};
    assign wire569 = {5'd4, 5'd2};
    assign wire570 = {5'd4, 5'd2};
    assign wire571 = {5'd4, 5'd2};
    assign wire572 = {5'd4, 5'd2};
    assign wire573 = {5'd4, 5'd2};
    assign wire574 = {5'd4, 5'd2};
    assign wire575 = {5'd4, 5'd2};
    assign wire576 = {5'd6, 5'd2};
    assign wire577 = {5'd6, 5'd2};
    assign wire578 = {5'd6, 5'd2};
    assign wire579 = {5'd6, 5'd2};
    assign wire580 = {5'd6, 5'd2};
    assign wire581 = {5'd6, 5'd2};
    assign wire582 = {5'd6, 5'd2};
    assign wire583 = {5'd6, 5'd2};
    assign wire584 = {5'd6, 5'd2};
    assign wire585 = {5'd6, 5'd2};
    assign wire586 = {5'd6, 5'd2};
    assign wire587 = {5'd6, 5'd2};
    assign wire588 = {5'd6, 5'd2};
    assign wire589 = {5'd6, 5'd2};
    assign wire590 = {5'd6, 5'd2};
    assign wire591 = {5'd6, 5'd2};
    assign wire592 = {5'd6, 5'd2};
    assign wire593 = {5'd6, 5'd2};
    assign wire594 = {5'd6, 5'd2};
    assign wire595 = {5'd6, 5'd2};
    assign wire596 = {5'd6, 5'd2};
    assign wire597 = {5'd6, 5'd2};
    assign wire598 = {5'd6, 5'd2};
    assign wire599 = {5'd6, 5'd2};
    assign wire600 = {5'd6, 5'd2};
    assign wire601 = {5'd6, 5'd2};
    assign wire602 = {5'd6, 5'd2};
    assign wire603 = {5'd6, 5'd2};
    assign wire604 = {5'd6, 5'd2};
    assign wire605 = {5'd6, 5'd2};
    assign wire606 = {5'd6, 5'd2};
    assign wire607 = {5'd6, 5'd2};
    assign wire608 = {5'd8, 5'd2};
    assign wire609 = {5'd8, 5'd2};
    assign wire610 = {5'd8, 5'd2};
    assign wire611 = {5'd8, 5'd2};
    assign wire612 = {5'd8, 5'd2};
    assign wire613 = {5'd8, 5'd2};
    assign wire614 = {5'd8, 5'd2};
    assign wire615 = {5'd8, 5'd2};
    assign wire616 = {5'd8, 5'd2};
    assign wire617 = {5'd8, 5'd2};
    assign wire618 = {5'd8, 5'd2};
    assign wire619 = {5'd8, 5'd2};
    assign wire620 = {5'd8, 5'd2};
    assign wire621 = {5'd8, 5'd2};
    assign wire622 = {5'd8, 5'd2};
    assign wire623 = {5'd8, 5'd2};
    assign wire624 = {5'd8, 5'd2};
    assign wire625 = {5'd8, 5'd2};
    assign wire626 = {5'd8, 5'd2};
    assign wire627 = {5'd8, 5'd2};
    assign wire628 = {5'd8, 5'd2};
    assign wire629 = {5'd8, 5'd2};
    assign wire630 = {5'd8, 5'd2};
    assign wire631 = {5'd8, 5'd2};
    assign wire632 = {5'd8, 5'd2};
    assign wire633 = {5'd8, 5'd2};
    assign wire634 = {5'd8, 5'd2};
    assign wire635 = {5'd8, 5'd2};
    assign wire636 = {5'd8, 5'd2};
    assign wire637 = {5'd8, 5'd2};
    assign wire638 = {5'd8, 5'd2};
    assign wire639 = {5'd8, 5'd2};
    assign wire640 = {5'd4, 5'd3};
    assign wire641 = {5'd4, 5'd3};
    assign wire642 = {5'd4, 5'd3};
    assign wire643 = {5'd4, 5'd3};
    assign wire644 = {5'd4, 5'd3};
    assign wire645 = {5'd6, 5'd5};
    assign wire646 = {5'd4, 5'd3};
    assign wire647 = {5'd4, 5'd3};
    assign wire648 = {5'd5, 5'd4};
    assign wire649 = {5'd5, 5'd4};
    assign wire650 = {5'd5, 5'd4};
    assign wire651 = {5'd5, 5'd4};
    assign wire652 = {5'd5, 5'd4};
    assign wire653 = {5'd5, 5'd4};
    assign wire654 = {5'd5, 5'd4};
    assign wire655 = {5'd5, 5'd4};
    assign wire656 = {5'd6, 5'd5};
    assign wire657 = {5'd6, 5'd5};
    assign wire658 = {5'd6, 5'd5};
    assign wire659 = {5'd6, 5'd5};
    assign wire660 = {5'd6, 5'd5};
    assign wire661 = {5'd6, 5'd5};
    assign wire662 = {5'd6, 5'd5};
    assign wire663 = {5'd6, 5'd5};
    assign wire664 = {5'd4, 5'd3};
    assign wire665 = {5'd4, 5'd3};
    assign wire666 = {5'd4, 5'd3};
    assign wire667 = {5'd4, 5'd3};
    assign wire668 = {5'd4, 5'd3};
    assign wire669 = {5'd4, 5'd3};
    assign wire670 = {5'd4, 5'd3};
    assign wire671 = {5'd4, 5'd3};
    assign wire672 = {5'd5, 5'd3};
    assign wire673 = {5'd5, 5'd3};
    assign wire674 = {5'd5, 5'd3};
    assign wire675 = {5'd5, 5'd3};
    assign wire676 = {5'd5, 5'd3};
    assign wire677 = {5'd7, 5'd5};
    assign wire678 = {5'd5, 5'd3};
    assign wire679 = {5'd5, 5'd3};
    assign wire680 = {5'd6, 5'd4};
    assign wire681 = {5'd6, 5'd4};
    assign wire682 = {5'd6, 5'd4};
    assign wire683 = {5'd6, 5'd4};
    assign wire684 = {5'd6, 5'd4};
    assign wire685 = {5'd6, 5'd4};
    assign wire686 = {5'd6, 5'd4};
    assign wire687 = {5'd6, 5'd4};
    assign wire688 = {5'd7, 5'd5};
    assign wire689 = {5'd7, 5'd5};
    assign wire690 = {5'd7, 5'd5};
    assign wire691 = {5'd7, 5'd5};
    assign wire692 = {5'd7, 5'd5};
    assign wire693 = {5'd7, 5'd5};
    assign wire694 = {5'd7, 5'd5};
    assign wire695 = {5'd7, 5'd5};
    assign wire696 = {5'd5, 5'd3};
    assign wire697 = {5'd5, 5'd3};
    assign wire698 = {5'd5, 5'd3};
    assign wire699 = {5'd5, 5'd3};
    assign wire700 = {5'd5, 5'd3};
    assign wire701 = {5'd5, 5'd3};
    assign wire702 = {5'd5, 5'd3};
    assign wire703 = {5'd5, 5'd3};
    assign wire704 = {5'd7, 5'd3};
    assign wire705 = {5'd7, 5'd3};
    assign wire706 = {5'd7, 5'd3};
    assign wire707 = {5'd7, 5'd3};
    assign wire708 = {5'd7, 5'd3};
    assign wire709 = {5'd9, 5'd5};
    assign wire710 = {5'd7, 5'd3};
    assign wire711 = {5'd7, 5'd3};
    assign wire712 = {5'd8, 5'd4};
    assign wire713 = {5'd8, 5'd4};
    assign wire714 = {5'd8, 5'd4};
    assign wire715 = {5'd8, 5'd4};
    assign wire716 = {5'd8, 5'd4};
    assign wire717 = {5'd8, 5'd4};
    assign wire718 = {5'd8, 5'd4};
    assign wire719 = {5'd8, 5'd4};
    assign wire720 = {5'd9, 5'd5};
    assign wire721 = {5'd9, 5'd5};
    assign wire722 = {5'd9, 5'd5};
    assign wire723 = {5'd9, 5'd5};
    assign wire724 = {5'd9, 5'd5};
    assign wire725 = {5'd9, 5'd5};
    assign wire726 = {5'd9, 5'd5};
    assign wire727 = {5'd9, 5'd5};
    assign wire728 = {5'd7, 5'd3};
    assign wire729 = {5'd7, 5'd3};
    assign wire730 = {5'd7, 5'd3};
    assign wire731 = {5'd7, 5'd3};
    assign wire732 = {5'd7, 5'd3};
    assign wire733 = {5'd7, 5'd3};
    assign wire734 = {5'd7, 5'd3};
    assign wire735 = {5'd7, 5'd3};
    assign wire736 = {5'd9, 5'd3};
    assign wire737 = {5'd9, 5'd3};
    assign wire738 = {5'd9, 5'd3};
    assign wire739 = {5'd9, 5'd3};
    assign wire740 = {5'd9, 5'd3};
    assign wire741 = {5'd11, 5'd5};
    assign wire742 = {5'd9, 5'd3};
    assign wire743 = {5'd9, 5'd3};
    assign wire744 = {5'd10, 5'd4};
    assign wire745 = {5'd10, 5'd4};
    assign wire746 = {5'd10, 5'd4};
    assign wire747 = {5'd10, 5'd4};
    assign wire748 = {5'd10, 5'd4};
    assign wire749 = {5'd10, 5'd4};
    assign wire750 = {5'd10, 5'd4};
    assign wire751 = {5'd10, 5'd4};
    assign wire752 = {5'd11, 5'd5};
    assign wire753 = {5'd11, 5'd5};
    assign wire754 = {5'd11, 5'd5};
    assign wire755 = {5'd11, 5'd5};
    assign wire756 = {5'd11, 5'd5};
    assign wire757 = {5'd11, 5'd5};
    assign wire758 = {5'd11, 5'd5};
    assign wire759 = {5'd11, 5'd5};
    assign wire760 = {5'd9, 5'd3};
    assign wire761 = {5'd9, 5'd3};
    assign wire762 = {5'd9, 5'd3};
    assign wire763 = {5'd9, 5'd3};
    assign wire764 = {5'd9, 5'd3};
    assign wire765 = {5'd9, 5'd3};
    assign wire766 = {5'd9, 5'd3};
    assign wire767 = {5'd9, 5'd3};
    assign wire768 = {5'd4, 5'd3};
    assign wire769 = {5'd4, 5'd3};
    assign wire770 = {5'd4, 5'd3};
    assign wire771 = {5'd4, 5'd3};
    assign wire772 = {5'd4, 5'd3};
    assign wire773 = {5'd4, 5'd3};
    assign wire774 = {5'd4, 5'd3};
    assign wire775 = {5'd4, 5'd3};
    assign wire776 = {5'd4, 5'd3};
    assign wire777 = {5'd4, 5'd3};
    assign wire778 = {5'd4, 5'd3};
    assign wire779 = {5'd4, 5'd3};
    assign wire780 = {5'd4, 5'd3};
    assign wire781 = {5'd4, 5'd3};
    assign wire782 = {5'd4, 5'd3};
    assign wire783 = {5'd4, 5'd3};
    assign wire784 = {5'd4, 5'd3};
    assign wire785 = {5'd4, 5'd3};
    assign wire786 = {5'd4, 5'd3};
    assign wire787 = {5'd4, 5'd3};
    assign wire788 = {5'd4, 5'd3};
    assign wire789 = {5'd4, 5'd3};
    assign wire790 = {5'd4, 5'd3};
    assign wire791 = {5'd4, 5'd3};
    assign wire792 = {5'd4, 5'd3};
    assign wire793 = {5'd4, 5'd3};
    assign wire794 = {5'd4, 5'd3};
    assign wire795 = {5'd4, 5'd3};
    assign wire796 = {5'd4, 5'd3};
    assign wire797 = {5'd4, 5'd3};
    assign wire798 = {5'd4, 5'd3};
    assign wire799 = {5'd4, 5'd3};
    assign wire800 = {5'd5, 5'd3};
    assign wire801 = {5'd5, 5'd3};
    assign wire802 = {5'd5, 5'd3};
    assign wire803 = {5'd5, 5'd3};
    assign wire804 = {5'd5, 5'd3};
    assign wire805 = {5'd5, 5'd3};
    assign wire806 = {5'd5, 5'd3};
    assign wire807 = {5'd5, 5'd3};
    assign wire808 = {5'd5, 5'd3};
    assign wire809 = {5'd5, 5'd3};
    assign wire810 = {5'd5, 5'd3};
    assign wire811 = {5'd5, 5'd3};
    assign wire812 = {5'd5, 5'd3};
    assign wire813 = {5'd5, 5'd3};
    assign wire814 = {5'd5, 5'd3};
    assign wire815 = {5'd5, 5'd3};
    assign wire816 = {5'd5, 5'd3};
    assign wire817 = {5'd5, 5'd3};
    assign wire818 = {5'd5, 5'd3};
    assign wire819 = {5'd5, 5'd3};
    assign wire820 = {5'd5, 5'd3};
    assign wire821 = {5'd5, 5'd3};
    assign wire822 = {5'd5, 5'd3};
    assign wire823 = {5'd5, 5'd3};
    assign wire824 = {5'd5, 5'd3};
    assign wire825 = {5'd5, 5'd3};
    assign wire826 = {5'd5, 5'd3};
    assign wire827 = {5'd5, 5'd3};
    assign wire828 = {5'd5, 5'd3};
    assign wire829 = {5'd5, 5'd3};
    assign wire830 = {5'd5, 5'd3};
    assign wire831 = {5'd5, 5'd3};
    assign wire832 = {5'd7, 5'd3};
    assign wire833 = {5'd7, 5'd3};
    assign wire834 = {5'd7, 5'd3};
    assign wire835 = {5'd7, 5'd3};
    assign wire836 = {5'd7, 5'd3};
    assign wire837 = {5'd7, 5'd3};
    assign wire838 = {5'd7, 5'd3};
    assign wire839 = {5'd7, 5'd3};
    assign wire840 = {5'd7, 5'd3};
    assign wire841 = {5'd7, 5'd3};
    assign wire842 = {5'd7, 5'd3};
    assign wire843 = {5'd7, 5'd3};
    assign wire844 = {5'd7, 5'd3};
    assign wire845 = {5'd7, 5'd3};
    assign wire846 = {5'd7, 5'd3};
    assign wire847 = {5'd7, 5'd3};
    assign wire848 = {5'd7, 5'd3};
    assign wire849 = {5'd7, 5'd3};
    assign wire850 = {5'd7, 5'd3};
    assign wire851 = {5'd7, 5'd3};
    assign wire852 = {5'd7, 5'd3};
    assign wire853 = {5'd7, 5'd3};
    assign wire854 = {5'd7, 5'd3};
    assign wire855 = {5'd7, 5'd3};
    assign wire856 = {5'd7, 5'd3};
    assign wire857 = {5'd7, 5'd3};
    assign wire858 = {5'd7, 5'd3};
    assign wire859 = {5'd7, 5'd3};
    assign wire860 = {5'd7, 5'd3};
    assign wire861 = {5'd7, 5'd3};
    assign wire862 = {5'd7, 5'd3};
    assign wire863 = {5'd7, 5'd3};
    assign wire864 = {5'd9, 5'd3};
    assign wire865 = {5'd9, 5'd3};
    assign wire866 = {5'd9, 5'd3};
    assign wire867 = {5'd9, 5'd3};
    assign wire868 = {5'd9, 5'd3};
    assign wire869 = {5'd9, 5'd3};
    assign wire870 = {5'd9, 5'd3};
    assign wire871 = {5'd9, 5'd3};
    assign wire872 = {5'd9, 5'd3};
    assign wire873 = {5'd9, 5'd3};
    assign wire874 = {5'd9, 5'd3};
    assign wire875 = {5'd9, 5'd3};
    assign wire876 = {5'd9, 5'd3};
    assign wire877 = {5'd9, 5'd3};
    assign wire878 = {5'd9, 5'd3};
    assign wire879 = {5'd9, 5'd3};
    assign wire880 = {5'd9, 5'd3};
    assign wire881 = {5'd9, 5'd3};
    assign wire882 = {5'd9, 5'd3};
    assign wire883 = {5'd9, 5'd3};
    assign wire884 = {5'd9, 5'd3};
    assign wire885 = {5'd9, 5'd3};
    assign wire886 = {5'd9, 5'd3};
    assign wire887 = {5'd9, 5'd3};
    assign wire888 = {5'd9, 5'd3};
    assign wire889 = {5'd9, 5'd3};
    assign wire890 = {5'd9, 5'd3};
    assign wire891 = {5'd9, 5'd3};
    assign wire892 = {5'd9, 5'd3};
    assign wire893 = {5'd9, 5'd3};
    assign wire894 = {5'd9, 5'd3};
    assign wire895 = {5'd9, 5'd3};
    assign wire896 = {5'd5, 5'd4};
    assign wire897 = {5'd5, 5'd4};
    assign wire898 = {5'd5, 5'd4};
    assign wire899 = {5'd5, 5'd4};
    assign wire900 = {5'd5, 5'd4};
    assign wire901 = {5'd7, 5'd6};
    assign wire902 = {5'd5, 5'd4};
    assign wire903 = {5'd5, 5'd4};
    assign wire904 = {5'd6, 5'd5};
    assign wire905 = {5'd6, 5'd5};
    assign wire906 = {5'd6, 5'd5};
    assign wire907 = {5'd6, 5'd5};
    assign wire908 = {5'd6, 5'd5};
    assign wire909 = {5'd6, 5'd5};
    assign wire910 = {5'd6, 5'd5};
    assign wire911 = {5'd6, 5'd5};
    assign wire912 = {5'd7, 5'd6};
    assign wire913 = {5'd7, 5'd6};
    assign wire914 = {5'd7, 5'd6};
    assign wire915 = {5'd7, 5'd6};
    assign wire916 = {5'd7, 5'd6};
    assign wire917 = {5'd7, 5'd6};
    assign wire918 = {5'd7, 5'd6};
    assign wire919 = {5'd7, 5'd6};
    assign wire920 = {5'd5, 5'd4};
    assign wire921 = {5'd5, 5'd4};
    assign wire922 = {5'd5, 5'd4};
    assign wire923 = {5'd5, 5'd4};
    assign wire924 = {5'd5, 5'd4};
    assign wire925 = {5'd5, 5'd4};
    assign wire926 = {5'd5, 5'd4};
    assign wire927 = {5'd5, 5'd4};
    assign wire928 = {5'd6, 5'd4};
    assign wire929 = {5'd6, 5'd4};
    assign wire930 = {5'd6, 5'd4};
    assign wire931 = {5'd6, 5'd4};
    assign wire932 = {5'd6, 5'd4};
    assign wire933 = {5'd8, 5'd6};
    assign wire934 = {5'd6, 5'd4};
    assign wire935 = {5'd6, 5'd4};
    assign wire936 = {5'd7, 5'd5};
    assign wire937 = {5'd7, 5'd5};
    assign wire938 = {5'd7, 5'd5};
    assign wire939 = {5'd7, 5'd5};
    assign wire940 = {5'd7, 5'd5};
    assign wire941 = {5'd7, 5'd5};
    assign wire942 = {5'd7, 5'd5};
    assign wire943 = {5'd7, 5'd5};
    assign wire944 = {5'd8, 5'd6};
    assign wire945 = {5'd8, 5'd6};
    assign wire946 = {5'd8, 5'd6};
    assign wire947 = {5'd8, 5'd6};
    assign wire948 = {5'd8, 5'd6};
    assign wire949 = {5'd8, 5'd6};
    assign wire950 = {5'd8, 5'd6};
    assign wire951 = {5'd8, 5'd6};
    assign wire952 = {5'd6, 5'd4};
    assign wire953 = {5'd6, 5'd4};
    assign wire954 = {5'd6, 5'd4};
    assign wire955 = {5'd6, 5'd4};
    assign wire956 = {5'd6, 5'd4};
    assign wire957 = {5'd6, 5'd4};
    assign wire958 = {5'd6, 5'd4};
    assign wire959 = {5'd6, 5'd4};
    assign wire960 = {5'd8, 5'd4};
    assign wire961 = {5'd8, 5'd4};
    assign wire962 = {5'd8, 5'd4};
    assign wire963 = {5'd8, 5'd4};
    assign wire964 = {5'd8, 5'd4};
    assign wire965 = {5'd10, 5'd6};
    assign wire966 = {5'd8, 5'd4};
    assign wire967 = {5'd8, 5'd4};
    assign wire968 = {5'd9, 5'd5};
    assign wire969 = {5'd9, 5'd5};
    assign wire970 = {5'd9, 5'd5};
    assign wire971 = {5'd9, 5'd5};
    assign wire972 = {5'd9, 5'd5};
    assign wire973 = {5'd9, 5'd5};
    assign wire974 = {5'd9, 5'd5};
    assign wire975 = {5'd9, 5'd5};
    assign wire976 = {5'd10, 5'd6};
    assign wire977 = {5'd10, 5'd6};
    assign wire978 = {5'd10, 5'd6};
    assign wire979 = {5'd10, 5'd6};
    assign wire980 = {5'd10, 5'd6};
    assign wire981 = {5'd10, 5'd6};
    assign wire982 = {5'd10, 5'd6};
    assign wire983 = {5'd10, 5'd6};
    assign wire984 = {5'd8, 5'd4};
    assign wire985 = {5'd8, 5'd4};
    assign wire986 = {5'd8, 5'd4};
    assign wire987 = {5'd8, 5'd4};
    assign wire988 = {5'd8, 5'd4};
    assign wire989 = {5'd8, 5'd4};
    assign wire990 = {5'd8, 5'd4};
    assign wire991 = {5'd8, 5'd4};
    assign wire992 = {5'd10, 5'd4};
    assign wire993 = {5'd10, 5'd4};
    assign wire994 = {5'd10, 5'd4};
    assign wire995 = {5'd10, 5'd4};
    assign wire996 = {5'd10, 5'd4};
    assign wire997 = {5'd12, 5'd6};
    assign wire998 = {5'd10, 5'd4};
    assign wire999 = {5'd10, 5'd4};
    assign wire1000 = {5'd11, 5'd5};
    assign wire1001 = {5'd11, 5'd5};
    assign wire1002 = {5'd11, 5'd5};
    assign wire1003 = {5'd11, 5'd5};
    assign wire1004 = {5'd11, 5'd5};
    assign wire1005 = {5'd11, 5'd5};
    assign wire1006 = {5'd11, 5'd5};
    assign wire1007 = {5'd11, 5'd5};
    assign wire1008 = {5'd12, 5'd6};
    assign wire1009 = {5'd12, 5'd6};
    assign wire1010 = {5'd12, 5'd6};
    assign wire1011 = {5'd12, 5'd6};
    assign wire1012 = {5'd12, 5'd6};
    assign wire1013 = {5'd12, 5'd6};
    assign wire1014 = {5'd12, 5'd6};
    assign wire1015 = {5'd12, 5'd6};
    assign wire1016 = {5'd10, 5'd4};
    assign wire1017 = {5'd10, 5'd4};
    assign wire1018 = {5'd10, 5'd4};
    assign wire1019 = {5'd10, 5'd4};
    assign wire1020 = {5'd10, 5'd4};
    assign wire1021 = {5'd10, 5'd4};
    assign wire1022 = {5'd10, 5'd4};
    assign wire1023 = {5'd10, 5'd4};
    assign wire1024 = {5'd3, 5'd2};
    assign wire1025 = {5'd3, 5'd2};
    assign wire1026 = {5'd3, 5'd2};
    assign wire1027 = {5'd3, 5'd2};
    assign wire1028 = {5'd3, 5'd2};
    assign wire1029 = {5'd3, 5'd2};
    assign wire1030 = {5'd3, 5'd2};
    assign wire1031 = {5'd3, 5'd2};
    assign wire1032 = {5'd3, 5'd2};
    assign wire1033 = {5'd3, 5'd2};
    assign wire1034 = {5'd3, 5'd2};
    assign wire1035 = {5'd3, 5'd2};
    assign wire1036 = {5'd3, 5'd2};
    assign wire1037 = {5'd3, 5'd2};
    assign wire1038 = {5'd3, 5'd2};
    assign wire1039 = {5'd3, 5'd2};
    assign wire1040 = {5'd3, 5'd2};
    assign wire1041 = {5'd3, 5'd2};
    assign wire1042 = {5'd3, 5'd2};
    assign wire1043 = {5'd3, 5'd2};
    assign wire1044 = {5'd3, 5'd2};
    assign wire1045 = {5'd3, 5'd2};
    assign wire1046 = {5'd3, 5'd2};
    assign wire1047 = {5'd3, 5'd2};
    assign wire1048 = {5'd3, 5'd2};
    assign wire1049 = {5'd3, 5'd2};
    assign wire1050 = {5'd3, 5'd2};
    assign wire1051 = {5'd3, 5'd2};
    assign wire1052 = {5'd3, 5'd2};
    assign wire1053 = {5'd3, 5'd2};
    assign wire1054 = {5'd3, 5'd2};
    assign wire1055 = {5'd3, 5'd2};
    assign wire1056 = {5'd4, 5'd2};
    assign wire1057 = {5'd4, 5'd2};
    assign wire1058 = {5'd4, 5'd2};
    assign wire1059 = {5'd4, 5'd2};
    assign wire1060 = {5'd4, 5'd2};
    assign wire1061 = {5'd4, 5'd2};
    assign wire1062 = {5'd4, 5'd2};
    assign wire1063 = {5'd4, 5'd2};
    assign wire1064 = {5'd4, 5'd2};
    assign wire1065 = {5'd4, 5'd2};
    assign wire1066 = {5'd4, 5'd2};
    assign wire1067 = {5'd4, 5'd2};
    assign wire1068 = {5'd4, 5'd2};
    assign wire1069 = {5'd4, 5'd2};
    assign wire1070 = {5'd4, 5'd2};
    assign wire1071 = {5'd4, 5'd2};
    assign wire1072 = {5'd4, 5'd2};
    assign wire1073 = {5'd4, 5'd2};
    assign wire1074 = {5'd4, 5'd2};
    assign wire1075 = {5'd4, 5'd2};
    assign wire1076 = {5'd4, 5'd2};
    assign wire1077 = {5'd4, 5'd2};
    assign wire1078 = {5'd4, 5'd2};
    assign wire1079 = {5'd4, 5'd2};
    assign wire1080 = {5'd4, 5'd2};
    assign wire1081 = {5'd4, 5'd2};
    assign wire1082 = {5'd4, 5'd2};
    assign wire1083 = {5'd4, 5'd2};
    assign wire1084 = {5'd4, 5'd2};
    assign wire1085 = {5'd4, 5'd2};
    assign wire1086 = {5'd4, 5'd2};
    assign wire1087 = {5'd4, 5'd2};
    assign wire1088 = {5'd6, 5'd2};
    assign wire1089 = {5'd6, 5'd2};
    assign wire1090 = {5'd6, 5'd2};
    assign wire1091 = {5'd6, 5'd2};
    assign wire1092 = {5'd6, 5'd2};
    assign wire1093 = {5'd6, 5'd2};
    assign wire1094 = {5'd6, 5'd2};
    assign wire1095 = {5'd6, 5'd2};
    assign wire1096 = {5'd6, 5'd2};
    assign wire1097 = {5'd6, 5'd2};
    assign wire1098 = {5'd6, 5'd2};
    assign wire1099 = {5'd6, 5'd2};
    assign wire1100 = {5'd6, 5'd2};
    assign wire1101 = {5'd6, 5'd2};
    assign wire1102 = {5'd6, 5'd2};
    assign wire1103 = {5'd6, 5'd2};
    assign wire1104 = {5'd6, 5'd2};
    assign wire1105 = {5'd6, 5'd2};
    assign wire1106 = {5'd6, 5'd2};
    assign wire1107 = {5'd6, 5'd2};
    assign wire1108 = {5'd6, 5'd2};
    assign wire1109 = {5'd6, 5'd2};
    assign wire1110 = {5'd6, 5'd2};
    assign wire1111 = {5'd6, 5'd2};
    assign wire1112 = {5'd6, 5'd2};
    assign wire1113 = {5'd6, 5'd2};
    assign wire1114 = {5'd6, 5'd2};
    assign wire1115 = {5'd6, 5'd2};
    assign wire1116 = {5'd6, 5'd2};
    assign wire1117 = {5'd6, 5'd2};
    assign wire1118 = {5'd6, 5'd2};
    assign wire1119 = {5'd6, 5'd2};
    assign wire1120 = {5'd8, 5'd2};
    assign wire1121 = {5'd8, 5'd2};
    assign wire1122 = {5'd8, 5'd2};
    assign wire1123 = {5'd8, 5'd2};
    assign wire1124 = {5'd8, 5'd2};
    assign wire1125 = {5'd8, 5'd2};
    assign wire1126 = {5'd8, 5'd2};
    assign wire1127 = {5'd8, 5'd2};
    assign wire1128 = {5'd8, 5'd2};
    assign wire1129 = {5'd8, 5'd2};
    assign wire1130 = {5'd8, 5'd2};
    assign wire1131 = {5'd8, 5'd2};
    assign wire1132 = {5'd8, 5'd2};
    assign wire1133 = {5'd8, 5'd2};
    assign wire1134 = {5'd8, 5'd2};
    assign wire1135 = {5'd8, 5'd2};
    assign wire1136 = {5'd8, 5'd2};
    assign wire1137 = {5'd8, 5'd2};
    assign wire1138 = {5'd8, 5'd2};
    assign wire1139 = {5'd8, 5'd2};
    assign wire1140 = {5'd8, 5'd2};
    assign wire1141 = {5'd8, 5'd2};
    assign wire1142 = {5'd8, 5'd2};
    assign wire1143 = {5'd8, 5'd2};
    assign wire1144 = {5'd8, 5'd2};
    assign wire1145 = {5'd8, 5'd2};
    assign wire1146 = {5'd8, 5'd2};
    assign wire1147 = {5'd8, 5'd2};
    assign wire1148 = {5'd8, 5'd2};
    assign wire1149 = {5'd8, 5'd2};
    assign wire1150 = {5'd8, 5'd2};
    assign wire1151 = {5'd8, 5'd2};
    assign wire1152 = {5'd4, 5'd3};
    assign wire1153 = {5'd4, 5'd3};
    assign wire1154 = {5'd4, 5'd3};
    assign wire1155 = {5'd4, 5'd3};
    assign wire1156 = {5'd5, 5'd4};
    assign wire1157 = {5'd8, 5'd7};
    assign wire1158 = {5'd4, 5'd3};
    assign wire1159 = {5'd4, 5'd3};
    assign wire1160 = {5'd5, 5'd4};
    assign wire1161 = {5'd5, 5'd4};
    assign wire1162 = {5'd5, 5'd4};
    assign wire1163 = {5'd5, 5'd4};
    assign wire1164 = {5'd6, 5'd5};
    assign wire1165 = {5'd5, 5'd4};
    assign wire1166 = {5'd5, 5'd4};
    assign wire1167 = {5'd5, 5'd4};
    assign wire1168 = {5'd8, 5'd7};
    assign wire1169 = {5'd8, 5'd7};
    assign wire1170 = {5'd8, 5'd7};
    assign wire1171 = {5'd8, 5'd7};
    assign wire1172 = {5'd9, 5'd8};
    assign wire1173 = {5'd8, 5'd7};
    assign wire1174 = {5'd8, 5'd7};
    assign wire1175 = {5'd8, 5'd7};
    assign wire1176 = {5'd4, 5'd3};
    assign wire1177 = {5'd4, 5'd3};
    assign wire1178 = {5'd4, 5'd3};
    assign wire1179 = {5'd4, 5'd3};
    assign wire1180 = {5'd4, 5'd3};
    assign wire1181 = {5'd4, 5'd3};
    assign wire1182 = {5'd4, 5'd3};
    assign wire1183 = {5'd4, 5'd3};
    assign wire1184 = {5'd5, 5'd3};
    assign wire1185 = {5'd5, 5'd3};
    assign wire1186 = {5'd5, 5'd3};
    assign wire1187 = {5'd5, 5'd3};
    assign wire1188 = {5'd6, 5'd4};
    assign wire1189 = {5'd9, 5'd7};
    assign wire1190 = {5'd5, 5'd3};
    assign wire1191 = {5'd5, 5'd3};
    assign wire1192 = {5'd6, 5'd4};
    assign wire1193 = {5'd6, 5'd4};
    assign wire1194 = {5'd6, 5'd4};
    assign wire1195 = {5'd6, 5'd4};
    assign wire1196 = {5'd7, 5'd5};
    assign wire1197 = {5'd6, 5'd4};
    assign wire1198 = {5'd6, 5'd4};
    assign wire1199 = {5'd6, 5'd4};
    assign wire1200 = {5'd9, 5'd7};
    assign wire1201 = {5'd9, 5'd7};
    assign wire1202 = {5'd9, 5'd7};
    assign wire1203 = {5'd9, 5'd7};
    assign wire1204 = {5'd10, 5'd8};
    assign wire1205 = {5'd9, 5'd7};
    assign wire1206 = {5'd9, 5'd7};
    assign wire1207 = {5'd9, 5'd7};
    assign wire1208 = {5'd5, 5'd3};
    assign wire1209 = {5'd5, 5'd3};
    assign wire1210 = {5'd5, 5'd3};
    assign wire1211 = {5'd5, 5'd3};
    assign wire1212 = {5'd5, 5'd3};
    assign wire1213 = {5'd5, 5'd3};
    assign wire1214 = {5'd5, 5'd3};
    assign wire1215 = {5'd5, 5'd3};
    assign wire1216 = {5'd7, 5'd3};
    assign wire1217 = {5'd7, 5'd3};
    assign wire1218 = {5'd7, 5'd3};
    assign wire1219 = {5'd7, 5'd3};
    assign wire1220 = {5'd8, 5'd4};
    assign wire1221 = {5'd11, 5'd7};
    assign wire1222 = {5'd7, 5'd3};
    assign wire1223 = {5'd7, 5'd3};
    assign wire1224 = {5'd8, 5'd4};
    assign wire1225 = {5'd8, 5'd4};
    assign wire1226 = {5'd8, 5'd4};
    assign wire1227 = {5'd8, 5'd4};
    assign wire1228 = {5'd9, 5'd5};
    assign wire1229 = {5'd8, 5'd4};
    assign wire1230 = {5'd8, 5'd4};
    assign wire1231 = {5'd8, 5'd4};
    assign wire1232 = {5'd11, 5'd7};
    assign wire1233 = {5'd11, 5'd7};
    assign wire1234 = {5'd11, 5'd7};
    assign wire1235 = {5'd11, 5'd7};
    assign wire1236 = {5'd12, 5'd8};
    assign wire1237 = {5'd11, 5'd7};
    assign wire1238 = {5'd11, 5'd7};
    assign wire1239 = {5'd11, 5'd7};
    assign wire1240 = {5'd7, 5'd3};
    assign wire1241 = {5'd7, 5'd3};
    assign wire1242 = {5'd7, 5'd3};
    assign wire1243 = {5'd7, 5'd3};
    assign wire1244 = {5'd7, 5'd3};
    assign wire1245 = {5'd7, 5'd3};
    assign wire1246 = {5'd7, 5'd3};
    assign wire1247 = {5'd7, 5'd3};
    assign wire1248 = {5'd9, 5'd3};
    assign wire1249 = {5'd9, 5'd3};
    assign wire1250 = {5'd9, 5'd3};
    assign wire1251 = {5'd9, 5'd3};
    assign wire1252 = {5'd10, 5'd4};
    assign wire1253 = {5'd13, 5'd7};
    assign wire1254 = {5'd9, 5'd3};
    assign wire1255 = {5'd9, 5'd3};
    assign wire1256 = {5'd10, 5'd4};
    assign wire1257 = {5'd10, 5'd4};
    assign wire1258 = {5'd10, 5'd4};
    assign wire1259 = {5'd10, 5'd4};
    assign wire1260 = {5'd11, 5'd5};
    assign wire1261 = {5'd10, 5'd4};
    assign wire1262 = {5'd10, 5'd4};
    assign wire1263 = {5'd10, 5'd4};
    assign wire1264 = {5'd13, 5'd7};
    assign wire1265 = {5'd13, 5'd7};
    assign wire1266 = {5'd13, 5'd7};
    assign wire1267 = {5'd13, 5'd7};
    assign wire1268 = {5'd14, 5'd8};
    assign wire1269 = {5'd13, 5'd7};
    assign wire1270 = {5'd13, 5'd7};
    assign wire1271 = {5'd13, 5'd7};
    assign wire1272 = {5'd9, 5'd3};
    assign wire1273 = {5'd9, 5'd3};
    assign wire1274 = {5'd9, 5'd3};
    assign wire1275 = {5'd9, 5'd3};
    assign wire1276 = {5'd9, 5'd3};
    assign wire1277 = {5'd9, 5'd3};
    assign wire1278 = {5'd9, 5'd3};
    assign wire1279 = {5'd9, 5'd3};
    assign wire1280 = {5'd4, 5'd3};
    assign wire1281 = {5'd4, 5'd3};
    assign wire1282 = {5'd4, 5'd3};
    assign wire1283 = {5'd4, 5'd3};
    assign wire1284 = {5'd4, 5'd3};
    assign wire1285 = {5'd4, 5'd3};
    assign wire1286 = {5'd4, 5'd3};
    assign wire1287 = {5'd4, 5'd3};
    assign wire1288 = {5'd4, 5'd3};
    assign wire1289 = {5'd4, 5'd3};
    assign wire1290 = {5'd4, 5'd3};
    assign wire1291 = {5'd4, 5'd3};
    assign wire1292 = {5'd4, 5'd3};
    assign wire1293 = {5'd4, 5'd3};
    assign wire1294 = {5'd4, 5'd3};
    assign wire1295 = {5'd4, 5'd3};
    assign wire1296 = {5'd4, 5'd3};
    assign wire1297 = {5'd4, 5'd3};
    assign wire1298 = {5'd4, 5'd3};
    assign wire1299 = {5'd4, 5'd3};
    assign wire1300 = {5'd4, 5'd3};
    assign wire1301 = {5'd4, 5'd3};
    assign wire1302 = {5'd4, 5'd3};
    assign wire1303 = {5'd4, 5'd3};
    assign wire1304 = {5'd4, 5'd3};
    assign wire1305 = {5'd4, 5'd3};
    assign wire1306 = {5'd4, 5'd3};
    assign wire1307 = {5'd4, 5'd3};
    assign wire1308 = {5'd4, 5'd3};
    assign wire1309 = {5'd4, 5'd3};
    assign wire1310 = {5'd4, 5'd3};
    assign wire1311 = {5'd4, 5'd3};
    assign wire1312 = {5'd5, 5'd3};
    assign wire1313 = {5'd5, 5'd3};
    assign wire1314 = {5'd5, 5'd3};
    assign wire1315 = {5'd5, 5'd3};
    assign wire1316 = {5'd5, 5'd3};
    assign wire1317 = {5'd5, 5'd3};
    assign wire1318 = {5'd5, 5'd3};
    assign wire1319 = {5'd5, 5'd3};
    assign wire1320 = {5'd5, 5'd3};
    assign wire1321 = {5'd5, 5'd3};
    assign wire1322 = {5'd5, 5'd3};
    assign wire1323 = {5'd5, 5'd3};
    assign wire1324 = {5'd5, 5'd3};
    assign wire1325 = {5'd5, 5'd3};
    assign wire1326 = {5'd5, 5'd3};
    assign wire1327 = {5'd5, 5'd3};
    assign wire1328 = {5'd5, 5'd3};
    assign wire1329 = {5'd5, 5'd3};
    assign wire1330 = {5'd5, 5'd3};
    assign wire1331 = {5'd5, 5'd3};
    assign wire1332 = {5'd5, 5'd3};
    assign wire1333 = {5'd5, 5'd3};
    assign wire1334 = {5'd5, 5'd3};
    assign wire1335 = {5'd5, 5'd3};
    assign wire1336 = {5'd5, 5'd3};
    assign wire1337 = {5'd5, 5'd3};
    assign wire1338 = {5'd5, 5'd3};
    assign wire1339 = {5'd5, 5'd3};
    assign wire1340 = {5'd5, 5'd3};
    assign wire1341 = {5'd5, 5'd3};
    assign wire1342 = {5'd5, 5'd3};
    assign wire1343 = {5'd5, 5'd3};
    assign wire1344 = {5'd7, 5'd3};
    assign wire1345 = {5'd7, 5'd3};
    assign wire1346 = {5'd7, 5'd3};
    assign wire1347 = {5'd7, 5'd3};
    assign wire1348 = {5'd7, 5'd3};
    assign wire1349 = {5'd7, 5'd3};
    assign wire1350 = {5'd7, 5'd3};
    assign wire1351 = {5'd7, 5'd3};
    assign wire1352 = {5'd7, 5'd3};
    assign wire1353 = {5'd7, 5'd3};
    assign wire1354 = {5'd7, 5'd3};
    assign wire1355 = {5'd7, 5'd3};
    assign wire1356 = {5'd7, 5'd3};
    assign wire1357 = {5'd7, 5'd3};
    assign wire1358 = {5'd7, 5'd3};
    assign wire1359 = {5'd7, 5'd3};
    assign wire1360 = {5'd7, 5'd3};
    assign wire1361 = {5'd7, 5'd3};
    assign wire1362 = {5'd7, 5'd3};
    assign wire1363 = {5'd7, 5'd3};
    assign wire1364 = {5'd7, 5'd3};
    assign wire1365 = {5'd7, 5'd3};
    assign wire1366 = {5'd7, 5'd3};
    assign wire1367 = {5'd7, 5'd3};
    assign wire1368 = {5'd7, 5'd3};
    assign wire1369 = {5'd7, 5'd3};
    assign wire1370 = {5'd7, 5'd3};
    assign wire1371 = {5'd7, 5'd3};
    assign wire1372 = {5'd7, 5'd3};
    assign wire1373 = {5'd7, 5'd3};
    assign wire1374 = {5'd7, 5'd3};
    assign wire1375 = {5'd7, 5'd3};
    assign wire1376 = {5'd9, 5'd3};
    assign wire1377 = {5'd9, 5'd3};
    assign wire1378 = {5'd9, 5'd3};
    assign wire1379 = {5'd9, 5'd3};
    assign wire1380 = {5'd9, 5'd3};
    assign wire1381 = {5'd9, 5'd3};
    assign wire1382 = {5'd9, 5'd3};
    assign wire1383 = {5'd9, 5'd3};
    assign wire1384 = {5'd9, 5'd3};
    assign wire1385 = {5'd9, 5'd3};
    assign wire1386 = {5'd9, 5'd3};
    assign wire1387 = {5'd9, 5'd3};
    assign wire1388 = {5'd9, 5'd3};
    assign wire1389 = {5'd9, 5'd3};
    assign wire1390 = {5'd9, 5'd3};
    assign wire1391 = {5'd9, 5'd3};
    assign wire1392 = {5'd9, 5'd3};
    assign wire1393 = {5'd9, 5'd3};
    assign wire1394 = {5'd9, 5'd3};
    assign wire1395 = {5'd9, 5'd3};
    assign wire1396 = {5'd9, 5'd3};
    assign wire1397 = {5'd9, 5'd3};
    assign wire1398 = {5'd9, 5'd3};
    assign wire1399 = {5'd9, 5'd3};
    assign wire1400 = {5'd9, 5'd3};
    assign wire1401 = {5'd9, 5'd3};
    assign wire1402 = {5'd9, 5'd3};
    assign wire1403 = {5'd9, 5'd3};
    assign wire1404 = {5'd9, 5'd3};
    assign wire1405 = {5'd9, 5'd3};
    assign wire1406 = {5'd9, 5'd3};
    assign wire1407 = {5'd9, 5'd3};
    assign wire1408 = {5'd5, 5'd4};
    assign wire1409 = {5'd5, 5'd4};
    assign wire1410 = {5'd5, 5'd4};
    assign wire1411 = {5'd5, 5'd4};
    assign wire1412 = {5'd6, 5'd5};
    assign wire1413 = {5'd9, 5'd8};
    assign wire1414 = {5'd5, 5'd4};
    assign wire1415 = {5'd5, 5'd4};
    assign wire1416 = {5'd6, 5'd5};
    assign wire1417 = {5'd6, 5'd5};
    assign wire1418 = {5'd6, 5'd5};
    assign wire1419 = {5'd6, 5'd5};
    assign wire1420 = {5'd7, 5'd6};
    assign wire1421 = {5'd6, 5'd5};
    assign wire1422 = {5'd6, 5'd5};
    assign wire1423 = {5'd6, 5'd5};
    assign wire1424 = {5'd9, 5'd8};
    assign wire1425 = {5'd9, 5'd8};
    assign wire1426 = {5'd9, 5'd8};
    assign wire1427 = {5'd9, 5'd8};
    assign wire1428 = {5'd10, 5'd9};
    assign wire1429 = {5'd9, 5'd8};
    assign wire1430 = {5'd9, 5'd8};
    assign wire1431 = {5'd9, 5'd8};
    assign wire1432 = {5'd5, 5'd4};
    assign wire1433 = {5'd5, 5'd4};
    assign wire1434 = {5'd5, 5'd4};
    assign wire1435 = {5'd5, 5'd4};
    assign wire1436 = {5'd5, 5'd4};
    assign wire1437 = {5'd5, 5'd4};
    assign wire1438 = {5'd5, 5'd4};
    assign wire1439 = {5'd5, 5'd4};
    assign wire1440 = {5'd6, 5'd4};
    assign wire1441 = {5'd6, 5'd4};
    assign wire1442 = {5'd6, 5'd4};
    assign wire1443 = {5'd6, 5'd4};
    assign wire1444 = {5'd7, 5'd5};
    assign wire1445 = {5'd10, 5'd8};
    assign wire1446 = {5'd6, 5'd4};
    assign wire1447 = {5'd6, 5'd4};
    assign wire1448 = {5'd7, 5'd5};
    assign wire1449 = {5'd7, 5'd5};
    assign wire1450 = {5'd7, 5'd5};
    assign wire1451 = {5'd7, 5'd5};
    assign wire1452 = {5'd8, 5'd6};
    assign wire1453 = {5'd7, 5'd5};
    assign wire1454 = {5'd7, 5'd5};
    assign wire1455 = {5'd7, 5'd5};
    assign wire1456 = {5'd10, 5'd8};
    assign wire1457 = {5'd10, 5'd8};
    assign wire1458 = {5'd10, 5'd8};
    assign wire1459 = {5'd10, 5'd8};
    assign wire1460 = {5'd11, 5'd9};
    assign wire1461 = {5'd10, 5'd8};
    assign wire1462 = {5'd10, 5'd8};
    assign wire1463 = {5'd10, 5'd8};
    assign wire1464 = {5'd6, 5'd4};
    assign wire1465 = {5'd6, 5'd4};
    assign wire1466 = {5'd6, 5'd4};
    assign wire1467 = {5'd6, 5'd4};
    assign wire1468 = {5'd6, 5'd4};
    assign wire1469 = {5'd6, 5'd4};
    assign wire1470 = {5'd6, 5'd4};
    assign wire1471 = {5'd6, 5'd4};
    assign wire1472 = {5'd8, 5'd4};
    assign wire1473 = {5'd8, 5'd4};
    assign wire1474 = {5'd8, 5'd4};
    assign wire1475 = {5'd8, 5'd4};
    assign wire1476 = {5'd9, 5'd5};
    assign wire1477 = {5'd12, 5'd8};
    assign wire1478 = {5'd8, 5'd4};
    assign wire1479 = {5'd8, 5'd4};
    assign wire1480 = {5'd9, 5'd5};
    assign wire1481 = {5'd9, 5'd5};
    assign wire1482 = {5'd9, 5'd5};
    assign wire1483 = {5'd9, 5'd5};
    assign wire1484 = {5'd10, 5'd6};
    assign wire1485 = {5'd9, 5'd5};
    assign wire1486 = {5'd9, 5'd5};
    assign wire1487 = {5'd9, 5'd5};
    assign wire1488 = {5'd12, 5'd8};
    assign wire1489 = {5'd12, 5'd8};
    assign wire1490 = {5'd12, 5'd8};
    assign wire1491 = {5'd12, 5'd8};
    assign wire1492 = {5'd13, 5'd9};
    assign wire1493 = {5'd12, 5'd8};
    assign wire1494 = {5'd12, 5'd8};
    assign wire1495 = {5'd12, 5'd8};
    assign wire1496 = {5'd8, 5'd4};
    assign wire1497 = {5'd8, 5'd4};
    assign wire1498 = {5'd8, 5'd4};
    assign wire1499 = {5'd8, 5'd4};
    assign wire1500 = {5'd8, 5'd4};
    assign wire1501 = {5'd8, 5'd4};
    assign wire1502 = {5'd8, 5'd4};
    assign wire1503 = {5'd8, 5'd4};
    assign wire1504 = {5'd10, 5'd4};
    assign wire1505 = {5'd10, 5'd4};
    assign wire1506 = {5'd10, 5'd4};
    assign wire1507 = {5'd10, 5'd4};
    assign wire1508 = {5'd11, 5'd5};
    assign wire1509 = {5'd14, 5'd8};
    assign wire1510 = {5'd10, 5'd4};
    assign wire1511 = {5'd10, 5'd4};
    assign wire1512 = {5'd11, 5'd5};
    assign wire1513 = {5'd11, 5'd5};
    assign wire1514 = {5'd11, 5'd5};
    assign wire1515 = {5'd11, 5'd5};
    assign wire1516 = {5'd12, 5'd6};
    assign wire1517 = {5'd11, 5'd5};
    assign wire1518 = {5'd11, 5'd5};
    assign wire1519 = {5'd11, 5'd5};
    assign wire1520 = {5'd14, 5'd8};
    assign wire1521 = {5'd14, 5'd8};
    assign wire1522 = {5'd14, 5'd8};
    assign wire1523 = {5'd14, 5'd8};
    assign wire1524 = {5'd15, 5'd9};
    assign wire1525 = {5'd14, 5'd8};
    assign wire1526 = {5'd14, 5'd8};
    assign wire1527 = {5'd14, 5'd8};
    assign wire1528 = {5'd10, 5'd4};
    assign wire1529 = {5'd10, 5'd4};
    assign wire1530 = {5'd10, 5'd4};
    assign wire1531 = {5'd10, 5'd4};
    assign wire1532 = {5'd10, 5'd4};
    assign wire1533 = {5'd10, 5'd4};
    assign wire1534 = {5'd10, 5'd4};
    assign wire1535 = {5'd10, 5'd4};
    assign wire1536 = {5'd4, 5'd3};
    assign wire1537 = {5'd4, 5'd3};
    assign wire1538 = {5'd4, 5'd3};
    assign wire1539 = {5'd4, 5'd3};
    assign wire1540 = {5'd4, 5'd3};
    assign wire1541 = {5'd4, 5'd3};
    assign wire1542 = {5'd4, 5'd3};
    assign wire1543 = {5'd4, 5'd3};
    assign wire1544 = {5'd4, 5'd3};
    assign wire1545 = {5'd4, 5'd3};
    assign wire1546 = {5'd4, 5'd3};
    assign wire1547 = {5'd4, 5'd3};
    assign wire1548 = {5'd4, 5'd3};
    assign wire1549 = {5'd4, 5'd3};
    assign wire1550 = {5'd4, 5'd3};
    assign wire1551 = {5'd4, 5'd3};
    assign wire1552 = {5'd4, 5'd3};
    assign wire1553 = {5'd4, 5'd3};
    assign wire1554 = {5'd4, 5'd3};
    assign wire1555 = {5'd4, 5'd3};
    assign wire1556 = {5'd4, 5'd3};
    assign wire1557 = {5'd4, 5'd3};
    assign wire1558 = {5'd4, 5'd3};
    assign wire1559 = {5'd4, 5'd3};
    assign wire1560 = {5'd4, 5'd3};
    assign wire1561 = {5'd4, 5'd3};
    assign wire1562 = {5'd4, 5'd3};
    assign wire1563 = {5'd4, 5'd3};
    assign wire1564 = {5'd4, 5'd3};
    assign wire1565 = {5'd4, 5'd3};
    assign wire1566 = {5'd4, 5'd3};
    assign wire1567 = {5'd4, 5'd3};
    assign wire1568 = {5'd5, 5'd3};
    assign wire1569 = {5'd5, 5'd3};
    assign wire1570 = {5'd5, 5'd3};
    assign wire1571 = {5'd5, 5'd3};
    assign wire1572 = {5'd5, 5'd3};
    assign wire1573 = {5'd5, 5'd3};
    assign wire1574 = {5'd5, 5'd3};
    assign wire1575 = {5'd5, 5'd3};
    assign wire1576 = {5'd5, 5'd3};
    assign wire1577 = {5'd5, 5'd3};
    assign wire1578 = {5'd5, 5'd3};
    assign wire1579 = {5'd5, 5'd3};
    assign wire1580 = {5'd5, 5'd3};
    assign wire1581 = {5'd5, 5'd3};
    assign wire1582 = {5'd5, 5'd3};
    assign wire1583 = {5'd5, 5'd3};
    assign wire1584 = {5'd5, 5'd3};
    assign wire1585 = {5'd5, 5'd3};
    assign wire1586 = {5'd5, 5'd3};
    assign wire1587 = {5'd5, 5'd3};
    assign wire1588 = {5'd5, 5'd3};
    assign wire1589 = {5'd5, 5'd3};
    assign wire1590 = {5'd5, 5'd3};
    assign wire1591 = {5'd5, 5'd3};
    assign wire1592 = {5'd5, 5'd3};
    assign wire1593 = {5'd5, 5'd3};
    assign wire1594 = {5'd5, 5'd3};
    assign wire1595 = {5'd5, 5'd3};
    assign wire1596 = {5'd5, 5'd3};
    assign wire1597 = {5'd5, 5'd3};
    assign wire1598 = {5'd5, 5'd3};
    assign wire1599 = {5'd5, 5'd3};
    assign wire1600 = {5'd7, 5'd3};
    assign wire1601 = {5'd7, 5'd3};
    assign wire1602 = {5'd7, 5'd3};
    assign wire1603 = {5'd7, 5'd3};
    assign wire1604 = {5'd7, 5'd3};
    assign wire1605 = {5'd7, 5'd3};
    assign wire1606 = {5'd7, 5'd3};
    assign wire1607 = {5'd7, 5'd3};
    assign wire1608 = {5'd7, 5'd3};
    assign wire1609 = {5'd7, 5'd3};
    assign wire1610 = {5'd7, 5'd3};
    assign wire1611 = {5'd7, 5'd3};
    assign wire1612 = {5'd7, 5'd3};
    assign wire1613 = {5'd7, 5'd3};
    assign wire1614 = {5'd7, 5'd3};
    assign wire1615 = {5'd7, 5'd3};
    assign wire1616 = {5'd7, 5'd3};
    assign wire1617 = {5'd7, 5'd3};
    assign wire1618 = {5'd7, 5'd3};
    assign wire1619 = {5'd7, 5'd3};
    assign wire1620 = {5'd7, 5'd3};
    assign wire1621 = {5'd7, 5'd3};
    assign wire1622 = {5'd7, 5'd3};
    assign wire1623 = {5'd7, 5'd3};
    assign wire1624 = {5'd7, 5'd3};
    assign wire1625 = {5'd7, 5'd3};
    assign wire1626 = {5'd7, 5'd3};
    assign wire1627 = {5'd7, 5'd3};
    assign wire1628 = {5'd7, 5'd3};
    assign wire1629 = {5'd7, 5'd3};
    assign wire1630 = {5'd7, 5'd3};
    assign wire1631 = {5'd7, 5'd3};
    assign wire1632 = {5'd9, 5'd3};
    assign wire1633 = {5'd9, 5'd3};
    assign wire1634 = {5'd9, 5'd3};
    assign wire1635 = {5'd9, 5'd3};
    assign wire1636 = {5'd9, 5'd3};
    assign wire1637 = {5'd9, 5'd3};
    assign wire1638 = {5'd9, 5'd3};
    assign wire1639 = {5'd9, 5'd3};
    assign wire1640 = {5'd9, 5'd3};
    assign wire1641 = {5'd9, 5'd3};
    assign wire1642 = {5'd9, 5'd3};
    assign wire1643 = {5'd9, 5'd3};
    assign wire1644 = {5'd9, 5'd3};
    assign wire1645 = {5'd9, 5'd3};
    assign wire1646 = {5'd9, 5'd3};
    assign wire1647 = {5'd9, 5'd3};
    assign wire1648 = {5'd9, 5'd3};
    assign wire1649 = {5'd9, 5'd3};
    assign wire1650 = {5'd9, 5'd3};
    assign wire1651 = {5'd9, 5'd3};
    assign wire1652 = {5'd9, 5'd3};
    assign wire1653 = {5'd9, 5'd3};
    assign wire1654 = {5'd9, 5'd3};
    assign wire1655 = {5'd9, 5'd3};
    assign wire1656 = {5'd9, 5'd3};
    assign wire1657 = {5'd9, 5'd3};
    assign wire1658 = {5'd9, 5'd3};
    assign wire1659 = {5'd9, 5'd3};
    assign wire1660 = {5'd9, 5'd3};
    assign wire1661 = {5'd9, 5'd3};
    assign wire1662 = {5'd9, 5'd3};
    assign wire1663 = {5'd9, 5'd3};
    assign wire1664 = {5'd5, 5'd4};
    assign wire1665 = {5'd5, 5'd4};
    assign wire1666 = {5'd5, 5'd4};
    assign wire1667 = {5'd5, 5'd4};
    assign wire1668 = {5'd5, 5'd4};
    assign wire1669 = {5'd7, 5'd6};
    assign wire1670 = {5'd5, 5'd4};
    assign wire1671 = {5'd5, 5'd4};
    assign wire1672 = {5'd6, 5'd5};
    assign wire1673 = {5'd6, 5'd5};
    assign wire1674 = {5'd6, 5'd5};
    assign wire1675 = {5'd6, 5'd5};
    assign wire1676 = {5'd6, 5'd5};
    assign wire1677 = {5'd6, 5'd5};
    assign wire1678 = {5'd6, 5'd5};
    assign wire1679 = {5'd6, 5'd5};
    assign wire1680 = {5'd7, 5'd6};
    assign wire1681 = {5'd7, 5'd6};
    assign wire1682 = {5'd7, 5'd6};
    assign wire1683 = {5'd7, 5'd6};
    assign wire1684 = {5'd7, 5'd6};
    assign wire1685 = {5'd7, 5'd6};
    assign wire1686 = {5'd7, 5'd6};
    assign wire1687 = {5'd7, 5'd6};
    assign wire1688 = {5'd5, 5'd4};
    assign wire1689 = {5'd5, 5'd4};
    assign wire1690 = {5'd5, 5'd4};
    assign wire1691 = {5'd5, 5'd4};
    assign wire1692 = {5'd5, 5'd4};
    assign wire1693 = {5'd5, 5'd4};
    assign wire1694 = {5'd5, 5'd4};
    assign wire1695 = {5'd5, 5'd4};
    assign wire1696 = {5'd6, 5'd4};
    assign wire1697 = {5'd6, 5'd4};
    assign wire1698 = {5'd6, 5'd4};
    assign wire1699 = {5'd6, 5'd4};
    assign wire1700 = {5'd6, 5'd4};
    assign wire1701 = {5'd8, 5'd6};
    assign wire1702 = {5'd6, 5'd4};
    assign wire1703 = {5'd6, 5'd4};
    assign wire1704 = {5'd7, 5'd5};
    assign wire1705 = {5'd7, 5'd5};
    assign wire1706 = {5'd7, 5'd5};
    assign wire1707 = {5'd7, 5'd5};
    assign wire1708 = {5'd7, 5'd5};
    assign wire1709 = {5'd7, 5'd5};
    assign wire1710 = {5'd7, 5'd5};
    assign wire1711 = {5'd7, 5'd5};
    assign wire1712 = {5'd8, 5'd6};
    assign wire1713 = {5'd8, 5'd6};
    assign wire1714 = {5'd8, 5'd6};
    assign wire1715 = {5'd8, 5'd6};
    assign wire1716 = {5'd8, 5'd6};
    assign wire1717 = {5'd8, 5'd6};
    assign wire1718 = {5'd8, 5'd6};
    assign wire1719 = {5'd8, 5'd6};
    assign wire1720 = {5'd6, 5'd4};
    assign wire1721 = {5'd6, 5'd4};
    assign wire1722 = {5'd6, 5'd4};
    assign wire1723 = {5'd6, 5'd4};
    assign wire1724 = {5'd6, 5'd4};
    assign wire1725 = {5'd6, 5'd4};
    assign wire1726 = {5'd6, 5'd4};
    assign wire1727 = {5'd6, 5'd4};
    assign wire1728 = {5'd8, 5'd4};
    assign wire1729 = {5'd8, 5'd4};
    assign wire1730 = {5'd8, 5'd4};
    assign wire1731 = {5'd8, 5'd4};
    assign wire1732 = {5'd8, 5'd4};
    assign wire1733 = {5'd10, 5'd6};
    assign wire1734 = {5'd8, 5'd4};
    assign wire1735 = {5'd8, 5'd4};
    assign wire1736 = {5'd9, 5'd5};
    assign wire1737 = {5'd9, 5'd5};
    assign wire1738 = {5'd9, 5'd5};
    assign wire1739 = {5'd9, 5'd5};
    assign wire1740 = {5'd9, 5'd5};
    assign wire1741 = {5'd9, 5'd5};
    assign wire1742 = {5'd9, 5'd5};
    assign wire1743 = {5'd9, 5'd5};
    assign wire1744 = {5'd10, 5'd6};
    assign wire1745 = {5'd10, 5'd6};
    assign wire1746 = {5'd10, 5'd6};
    assign wire1747 = {5'd10, 5'd6};
    assign wire1748 = {5'd10, 5'd6};
    assign wire1749 = {5'd10, 5'd6};
    assign wire1750 = {5'd10, 5'd6};
    assign wire1751 = {5'd10, 5'd6};
    assign wire1752 = {5'd8, 5'd4};
    assign wire1753 = {5'd8, 5'd4};
    assign wire1754 = {5'd8, 5'd4};
    assign wire1755 = {5'd8, 5'd4};
    assign wire1756 = {5'd8, 5'd4};
    assign wire1757 = {5'd8, 5'd4};
    assign wire1758 = {5'd8, 5'd4};
    assign wire1759 = {5'd8, 5'd4};
    assign wire1760 = {5'd10, 5'd4};
    assign wire1761 = {5'd10, 5'd4};
    assign wire1762 = {5'd10, 5'd4};
    assign wire1763 = {5'd10, 5'd4};
    assign wire1764 = {5'd10, 5'd4};
    assign wire1765 = {5'd12, 5'd6};
    assign wire1766 = {5'd10, 5'd4};
    assign wire1767 = {5'd10, 5'd4};
    assign wire1768 = {5'd11, 5'd5};
    assign wire1769 = {5'd11, 5'd5};
    assign wire1770 = {5'd11, 5'd5};
    assign wire1771 = {5'd11, 5'd5};
    assign wire1772 = {5'd11, 5'd5};
    assign wire1773 = {5'd11, 5'd5};
    assign wire1774 = {5'd11, 5'd5};
    assign wire1775 = {5'd11, 5'd5};
    assign wire1776 = {5'd12, 5'd6};
    assign wire1777 = {5'd12, 5'd6};
    assign wire1778 = {5'd12, 5'd6};
    assign wire1779 = {5'd12, 5'd6};
    assign wire1780 = {5'd12, 5'd6};
    assign wire1781 = {5'd12, 5'd6};
    assign wire1782 = {5'd12, 5'd6};
    assign wire1783 = {5'd12, 5'd6};
    assign wire1784 = {5'd10, 5'd4};
    assign wire1785 = {5'd10, 5'd4};
    assign wire1786 = {5'd10, 5'd4};
    assign wire1787 = {5'd10, 5'd4};
    assign wire1788 = {5'd10, 5'd4};
    assign wire1789 = {5'd10, 5'd4};
    assign wire1790 = {5'd10, 5'd4};
    assign wire1791 = {5'd10, 5'd4};
    assign wire1792 = {5'd5, 5'd4};
    assign wire1793 = {5'd5, 5'd4};
    assign wire1794 = {5'd5, 5'd4};
    assign wire1795 = {5'd5, 5'd4};
    assign wire1796 = {5'd5, 5'd4};
    assign wire1797 = {5'd5, 5'd4};
    assign wire1798 = {5'd5, 5'd4};
    assign wire1799 = {5'd5, 5'd4};
    assign wire1800 = {5'd5, 5'd4};
    assign wire1801 = {5'd5, 5'd4};
    assign wire1802 = {5'd5, 5'd4};
    assign wire1803 = {5'd5, 5'd4};
    assign wire1804 = {5'd5, 5'd4};
    assign wire1805 = {5'd5, 5'd4};
    assign wire1806 = {5'd5, 5'd4};
    assign wire1807 = {5'd5, 5'd4};
    assign wire1808 = {5'd5, 5'd4};
    assign wire1809 = {5'd5, 5'd4};
    assign wire1810 = {5'd5, 5'd4};
    assign wire1811 = {5'd5, 5'd4};
    assign wire1812 = {5'd5, 5'd4};
    assign wire1813 = {5'd5, 5'd4};
    assign wire1814 = {5'd5, 5'd4};
    assign wire1815 = {5'd5, 5'd4};
    assign wire1816 = {5'd5, 5'd4};
    assign wire1817 = {5'd5, 5'd4};
    assign wire1818 = {5'd5, 5'd4};
    assign wire1819 = {5'd5, 5'd4};
    assign wire1820 = {5'd5, 5'd4};
    assign wire1821 = {5'd5, 5'd4};
    assign wire1822 = {5'd5, 5'd4};
    assign wire1823 = {5'd5, 5'd4};
    assign wire1824 = {5'd6, 5'd4};
    assign wire1825 = {5'd6, 5'd4};
    assign wire1826 = {5'd6, 5'd4};
    assign wire1827 = {5'd6, 5'd4};
    assign wire1828 = {5'd6, 5'd4};
    assign wire1829 = {5'd6, 5'd4};
    assign wire1830 = {5'd6, 5'd4};
    assign wire1831 = {5'd6, 5'd4};
    assign wire1832 = {5'd6, 5'd4};
    assign wire1833 = {5'd6, 5'd4};
    assign wire1834 = {5'd6, 5'd4};
    assign wire1835 = {5'd6, 5'd4};
    assign wire1836 = {5'd6, 5'd4};
    assign wire1837 = {5'd6, 5'd4};
    assign wire1838 = {5'd6, 5'd4};
    assign wire1839 = {5'd6, 5'd4};
    assign wire1840 = {5'd6, 5'd4};
    assign wire1841 = {5'd6, 5'd4};
    assign wire1842 = {5'd6, 5'd4};
    assign wire1843 = {5'd6, 5'd4};
    assign wire1844 = {5'd6, 5'd4};
    assign wire1845 = {5'd6, 5'd4};
    assign wire1846 = {5'd6, 5'd4};
    assign wire1847 = {5'd6, 5'd4};
    assign wire1848 = {5'd6, 5'd4};
    assign wire1849 = {5'd6, 5'd4};
    assign wire1850 = {5'd6, 5'd4};
    assign wire1851 = {5'd6, 5'd4};
    assign wire1852 = {5'd6, 5'd4};
    assign wire1853 = {5'd6, 5'd4};
    assign wire1854 = {5'd6, 5'd4};
    assign wire1855 = {5'd6, 5'd4};
    assign wire1856 = {5'd8, 5'd4};
    assign wire1857 = {5'd8, 5'd4};
    assign wire1858 = {5'd8, 5'd4};
    assign wire1859 = {5'd8, 5'd4};
    assign wire1860 = {5'd8, 5'd4};
    assign wire1861 = {5'd8, 5'd4};
    assign wire1862 = {5'd8, 5'd4};
    assign wire1863 = {5'd8, 5'd4};
    assign wire1864 = {5'd8, 5'd4};
    assign wire1865 = {5'd8, 5'd4};
    assign wire1866 = {5'd8, 5'd4};
    assign wire1867 = {5'd8, 5'd4};
    assign wire1868 = {5'd8, 5'd4};
    assign wire1869 = {5'd8, 5'd4};
    assign wire1870 = {5'd8, 5'd4};
    assign wire1871 = {5'd8, 5'd4};
    assign wire1872 = {5'd8, 5'd4};
    assign wire1873 = {5'd8, 5'd4};
    assign wire1874 = {5'd8, 5'd4};
    assign wire1875 = {5'd8, 5'd4};
    assign wire1876 = {5'd8, 5'd4};
    assign wire1877 = {5'd8, 5'd4};
    assign wire1878 = {5'd8, 5'd4};
    assign wire1879 = {5'd8, 5'd4};
    assign wire1880 = {5'd8, 5'd4};
    assign wire1881 = {5'd8, 5'd4};
    assign wire1882 = {5'd8, 5'd4};
    assign wire1883 = {5'd8, 5'd4};
    assign wire1884 = {5'd8, 5'd4};
    assign wire1885 = {5'd8, 5'd4};
    assign wire1886 = {5'd8, 5'd4};
    assign wire1887 = {5'd8, 5'd4};
    assign wire1888 = {5'd10, 5'd4};
    assign wire1889 = {5'd10, 5'd4};
    assign wire1890 = {5'd10, 5'd4};
    assign wire1891 = {5'd10, 5'd4};
    assign wire1892 = {5'd10, 5'd4};
    assign wire1893 = {5'd10, 5'd4};
    assign wire1894 = {5'd10, 5'd4};
    assign wire1895 = {5'd10, 5'd4};
    assign wire1896 = {5'd10, 5'd4};
    assign wire1897 = {5'd10, 5'd4};
    assign wire1898 = {5'd10, 5'd4};
    assign wire1899 = {5'd10, 5'd4};
    assign wire1900 = {5'd10, 5'd4};
    assign wire1901 = {5'd10, 5'd4};
    assign wire1902 = {5'd10, 5'd4};
    assign wire1903 = {5'd10, 5'd4};
    assign wire1904 = {5'd10, 5'd4};
    assign wire1905 = {5'd10, 5'd4};
    assign wire1906 = {5'd10, 5'd4};
    assign wire1907 = {5'd10, 5'd4};
    assign wire1908 = {5'd10, 5'd4};
    assign wire1909 = {5'd10, 5'd4};
    assign wire1910 = {5'd10, 5'd4};
    assign wire1911 = {5'd10, 5'd4};
    assign wire1912 = {5'd10, 5'd4};
    assign wire1913 = {5'd10, 5'd4};
    assign wire1914 = {5'd10, 5'd4};
    assign wire1915 = {5'd10, 5'd4};
    assign wire1916 = {5'd10, 5'd4};
    assign wire1917 = {5'd10, 5'd4};
    assign wire1918 = {5'd10, 5'd4};
    assign wire1919 = {5'd10, 5'd4};
    assign wire1920 = {5'd6, 5'd5};
    assign wire1921 = {5'd6, 5'd5};
    assign wire1922 = {5'd6, 5'd5};
    assign wire1923 = {5'd6, 5'd5};
    assign wire1924 = {5'd6, 5'd5};
    assign wire1925 = {5'd8, 5'd7};
    assign wire1926 = {5'd6, 5'd5};
    assign wire1927 = {5'd6, 5'd5};
    assign wire1928 = {5'd7, 5'd6};
    assign wire1929 = {5'd7, 5'd6};
    assign wire1930 = {5'd7, 5'd6};
    assign wire1931 = {5'd7, 5'd6};
    assign wire1932 = {5'd7, 5'd6};
    assign wire1933 = {5'd7, 5'd6};
    assign wire1934 = {5'd7, 5'd6};
    assign wire1935 = {5'd7, 5'd6};
    assign wire1936 = {5'd8, 5'd7};
    assign wire1937 = {5'd8, 5'd7};
    assign wire1938 = {5'd8, 5'd7};
    assign wire1939 = {5'd8, 5'd7};
    assign wire1940 = {5'd8, 5'd7};
    assign wire1941 = {5'd8, 5'd7};
    assign wire1942 = {5'd8, 5'd7};
    assign wire1943 = {5'd8, 5'd7};
    assign wire1944 = {5'd6, 5'd5};
    assign wire1945 = {5'd6, 5'd5};
    assign wire1946 = {5'd6, 5'd5};
    assign wire1947 = {5'd6, 5'd5};
    assign wire1948 = {5'd6, 5'd5};
    assign wire1949 = {5'd6, 5'd5};
    assign wire1950 = {5'd6, 5'd5};
    assign wire1951 = {5'd6, 5'd5};
    assign wire1952 = {5'd7, 5'd5};
    assign wire1953 = {5'd7, 5'd5};
    assign wire1954 = {5'd7, 5'd5};
    assign wire1955 = {5'd7, 5'd5};
    assign wire1956 = {5'd7, 5'd5};
    assign wire1957 = {5'd9, 5'd7};
    assign wire1958 = {5'd7, 5'd5};
    assign wire1959 = {5'd7, 5'd5};
    assign wire1960 = {5'd8, 5'd6};
    assign wire1961 = {5'd8, 5'd6};
    assign wire1962 = {5'd8, 5'd6};
    assign wire1963 = {5'd8, 5'd6};
    assign wire1964 = {5'd8, 5'd6};
    assign wire1965 = {5'd8, 5'd6};
    assign wire1966 = {5'd8, 5'd6};
    assign wire1967 = {5'd8, 5'd6};
    assign wire1968 = {5'd9, 5'd7};
    assign wire1969 = {5'd9, 5'd7};
    assign wire1970 = {5'd9, 5'd7};
    assign wire1971 = {5'd9, 5'd7};
    assign wire1972 = {5'd9, 5'd7};
    assign wire1973 = {5'd9, 5'd7};
    assign wire1974 = {5'd9, 5'd7};
    assign wire1975 = {5'd9, 5'd7};
    assign wire1976 = {5'd7, 5'd5};
    assign wire1977 = {5'd7, 5'd5};
    assign wire1978 = {5'd7, 5'd5};
    assign wire1979 = {5'd7, 5'd5};
    assign wire1980 = {5'd7, 5'd5};
    assign wire1981 = {5'd7, 5'd5};
    assign wire1982 = {5'd7, 5'd5};
    assign wire1983 = {5'd7, 5'd5};
    assign wire1984 = {5'd9, 5'd5};
    assign wire1985 = {5'd9, 5'd5};
    assign wire1986 = {5'd9, 5'd5};
    assign wire1987 = {5'd9, 5'd5};
    assign wire1988 = {5'd9, 5'd5};
    assign wire1989 = {5'd11, 5'd7};
    assign wire1990 = {5'd9, 5'd5};
    assign wire1991 = {5'd9, 5'd5};
    assign wire1992 = {5'd10, 5'd6};
    assign wire1993 = {5'd10, 5'd6};
    assign wire1994 = {5'd10, 5'd6};
    assign wire1995 = {5'd10, 5'd6};
    assign wire1996 = {5'd10, 5'd6};
    assign wire1997 = {5'd10, 5'd6};
    assign wire1998 = {5'd10, 5'd6};
    assign wire1999 = {5'd10, 5'd6};
    assign wire2000 = {5'd11, 5'd7};
    assign wire2001 = {5'd11, 5'd7};
    assign wire2002 = {5'd11, 5'd7};
    assign wire2003 = {5'd11, 5'd7};
    assign wire2004 = {5'd11, 5'd7};
    assign wire2005 = {5'd11, 5'd7};
    assign wire2006 = {5'd11, 5'd7};
    assign wire2007 = {5'd11, 5'd7};
    assign wire2008 = {5'd9, 5'd5};
    assign wire2009 = {5'd9, 5'd5};
    assign wire2010 = {5'd9, 5'd5};
    assign wire2011 = {5'd9, 5'd5};
    assign wire2012 = {5'd9, 5'd5};
    assign wire2013 = {5'd9, 5'd5};
    assign wire2014 = {5'd9, 5'd5};
    assign wire2015 = {5'd9, 5'd5};
    assign wire2016 = {5'd11, 5'd5};
    assign wire2017 = {5'd11, 5'd5};
    assign wire2018 = {5'd11, 5'd5};
    assign wire2019 = {5'd11, 5'd5};
    assign wire2020 = {5'd11, 5'd5};
    assign wire2021 = {5'd13, 5'd7};
    assign wire2022 = {5'd11, 5'd5};
    assign wire2023 = {5'd11, 5'd5};
    assign wire2024 = {5'd12, 5'd6};
    assign wire2025 = {5'd12, 5'd6};
    assign wire2026 = {5'd12, 5'd6};
    assign wire2027 = {5'd12, 5'd6};
    assign wire2028 = {5'd12, 5'd6};
    assign wire2029 = {5'd12, 5'd6};
    assign wire2030 = {5'd12, 5'd6};
    assign wire2031 = {5'd12, 5'd6};
    assign wire2032 = {5'd13, 5'd7};
    assign wire2033 = {5'd13, 5'd7};
    assign wire2034 = {5'd13, 5'd7};
    assign wire2035 = {5'd13, 5'd7};
    assign wire2036 = {5'd13, 5'd7};
    assign wire2037 = {5'd13, 5'd7};
    assign wire2038 = {5'd13, 5'd7};
    assign wire2039 = {5'd13, 5'd7};
    assign wire2040 = {5'd11, 5'd5};
    assign wire2041 = {5'd11, 5'd5};
    assign wire2042 = {5'd11, 5'd5};
    assign wire2043 = {5'd11, 5'd5};
    assign wire2044 = {5'd11, 5'd5};
    assign wire2045 = {5'd11, 5'd5};
    assign wire2046 = {5'd11, 5'd5};
    assign wire2047 = {5'd11, 5'd5};
    assign wire2048 = {5'd3, 5'd2};
    assign wire2049 = {5'd3, 5'd2};
    assign wire2050 = {5'd3, 5'd2};
    assign wire2051 = {5'd3, 5'd2};
    assign wire2052 = {5'd3, 5'd2};
    assign wire2053 = {5'd3, 5'd2};
    assign wire2054 = {5'd3, 5'd2};
    assign wire2055 = {5'd3, 5'd2};
    assign wire2056 = {5'd3, 5'd2};
    assign wire2057 = {5'd3, 5'd2};
    assign wire2058 = {5'd3, 5'd2};
    assign wire2059 = {5'd3, 5'd2};
    assign wire2060 = {5'd3, 5'd2};
    assign wire2061 = {5'd3, 5'd2};
    assign wire2062 = {5'd3, 5'd2};
    assign wire2063 = {5'd3, 5'd2};
    assign wire2064 = {5'd3, 5'd2};
    assign wire2065 = {5'd3, 5'd2};
    assign wire2066 = {5'd3, 5'd2};
    assign wire2067 = {5'd3, 5'd2};
    assign wire2068 = {5'd3, 5'd2};
    assign wire2069 = {5'd3, 5'd2};
    assign wire2070 = {5'd3, 5'd2};
    assign wire2071 = {5'd3, 5'd2};
    assign wire2072 = {5'd3, 5'd2};
    assign wire2073 = {5'd3, 5'd2};
    assign wire2074 = {5'd3, 5'd2};
    assign wire2075 = {5'd3, 5'd2};
    assign wire2076 = {5'd3, 5'd2};
    assign wire2077 = {5'd3, 5'd2};
    assign wire2078 = {5'd3, 5'd2};
    assign wire2079 = {5'd3, 5'd2};
    assign wire2080 = {5'd4, 5'd2};
    assign wire2081 = {5'd4, 5'd2};
    assign wire2082 = {5'd4, 5'd2};
    assign wire2083 = {5'd4, 5'd2};
    assign wire2084 = {5'd4, 5'd2};
    assign wire2085 = {5'd4, 5'd2};
    assign wire2086 = {5'd4, 5'd2};
    assign wire2087 = {5'd4, 5'd2};
    assign wire2088 = {5'd4, 5'd2};
    assign wire2089 = {5'd4, 5'd2};
    assign wire2090 = {5'd4, 5'd2};
    assign wire2091 = {5'd4, 5'd2};
    assign wire2092 = {5'd4, 5'd2};
    assign wire2093 = {5'd4, 5'd2};
    assign wire2094 = {5'd4, 5'd2};
    assign wire2095 = {5'd4, 5'd2};
    assign wire2096 = {5'd4, 5'd2};
    assign wire2097 = {5'd4, 5'd2};
    assign wire2098 = {5'd4, 5'd2};
    assign wire2099 = {5'd4, 5'd2};
    assign wire2100 = {5'd4, 5'd2};
    assign wire2101 = {5'd4, 5'd2};
    assign wire2102 = {5'd4, 5'd2};
    assign wire2103 = {5'd4, 5'd2};
    assign wire2104 = {5'd4, 5'd2};
    assign wire2105 = {5'd4, 5'd2};
    assign wire2106 = {5'd4, 5'd2};
    assign wire2107 = {5'd4, 5'd2};
    assign wire2108 = {5'd4, 5'd2};
    assign wire2109 = {5'd4, 5'd2};
    assign wire2110 = {5'd4, 5'd2};
    assign wire2111 = {5'd4, 5'd2};
    assign wire2112 = {5'd6, 5'd2};
    assign wire2113 = {5'd6, 5'd2};
    assign wire2114 = {5'd6, 5'd2};
    assign wire2115 = {5'd6, 5'd2};
    assign wire2116 = {5'd6, 5'd2};
    assign wire2117 = {5'd6, 5'd2};
    assign wire2118 = {5'd6, 5'd2};
    assign wire2119 = {5'd6, 5'd2};
    assign wire2120 = {5'd6, 5'd2};
    assign wire2121 = {5'd6, 5'd2};
    assign wire2122 = {5'd6, 5'd2};
    assign wire2123 = {5'd6, 5'd2};
    assign wire2124 = {5'd6, 5'd2};
    assign wire2125 = {5'd6, 5'd2};
    assign wire2126 = {5'd6, 5'd2};
    assign wire2127 = {5'd6, 5'd2};
    assign wire2128 = {5'd6, 5'd2};
    assign wire2129 = {5'd6, 5'd2};
    assign wire2130 = {5'd6, 5'd2};
    assign wire2131 = {5'd6, 5'd2};
    assign wire2132 = {5'd6, 5'd2};
    assign wire2133 = {5'd6, 5'd2};
    assign wire2134 = {5'd6, 5'd2};
    assign wire2135 = {5'd6, 5'd2};
    assign wire2136 = {5'd6, 5'd2};
    assign wire2137 = {5'd6, 5'd2};
    assign wire2138 = {5'd6, 5'd2};
    assign wire2139 = {5'd6, 5'd2};
    assign wire2140 = {5'd6, 5'd2};
    assign wire2141 = {5'd6, 5'd2};
    assign wire2142 = {5'd6, 5'd2};
    assign wire2143 = {5'd6, 5'd2};
    assign wire2144 = {5'd8, 5'd2};
    assign wire2145 = {5'd8, 5'd2};
    assign wire2146 = {5'd8, 5'd2};
    assign wire2147 = {5'd8, 5'd2};
    assign wire2148 = {5'd8, 5'd2};
    assign wire2149 = {5'd8, 5'd2};
    assign wire2150 = {5'd8, 5'd2};
    assign wire2151 = {5'd8, 5'd2};
    assign wire2152 = {5'd8, 5'd2};
    assign wire2153 = {5'd8, 5'd2};
    assign wire2154 = {5'd8, 5'd2};
    assign wire2155 = {5'd8, 5'd2};
    assign wire2156 = {5'd8, 5'd2};
    assign wire2157 = {5'd8, 5'd2};
    assign wire2158 = {5'd8, 5'd2};
    assign wire2159 = {5'd8, 5'd2};
    assign wire2160 = {5'd8, 5'd2};
    assign wire2161 = {5'd8, 5'd2};
    assign wire2162 = {5'd8, 5'd2};
    assign wire2163 = {5'd8, 5'd2};
    assign wire2164 = {5'd8, 5'd2};
    assign wire2165 = {5'd8, 5'd2};
    assign wire2166 = {5'd8, 5'd2};
    assign wire2167 = {5'd8, 5'd2};
    assign wire2168 = {5'd8, 5'd2};
    assign wire2169 = {5'd8, 5'd2};
    assign wire2170 = {5'd8, 5'd2};
    assign wire2171 = {5'd8, 5'd2};
    assign wire2172 = {5'd8, 5'd2};
    assign wire2173 = {5'd8, 5'd2};
    assign wire2174 = {5'd8, 5'd2};
    assign wire2175 = {5'd8, 5'd2};
    assign wire2176 = {5'd4, 5'd3};
    assign wire2177 = {5'd4, 5'd3};
    assign wire2178 = {5'd4, 5'd3};
    assign wire2179 = {5'd4, 5'd3};
    assign wire2180 = {5'd5, 5'd4};
    assign wire2181 = {5'd8, 5'd7};
    assign wire2182 = {5'd4, 5'd3};
    assign wire2183 = {5'd4, 5'd3};
    assign wire2184 = {5'd5, 5'd4};
    assign wire2185 = {5'd5, 5'd4};
    assign wire2186 = {5'd5, 5'd4};
    assign wire2187 = {5'd5, 5'd4};
    assign wire2188 = {5'd6, 5'd5};
    assign wire2189 = {5'd5, 5'd4};
    assign wire2190 = {5'd5, 5'd4};
    assign wire2191 = {5'd5, 5'd4};
    assign wire2192 = {5'd8, 5'd7};
    assign wire2193 = {5'd8, 5'd7};
    assign wire2194 = {5'd8, 5'd7};
    assign wire2195 = {5'd8, 5'd7};
    assign wire2196 = {5'd9, 5'd8};
    assign wire2197 = {5'd8, 5'd7};
    assign wire2198 = {5'd8, 5'd7};
    assign wire2199 = {5'd8, 5'd7};
    assign wire2200 = {5'd4, 5'd3};
    assign wire2201 = {5'd4, 5'd3};
    assign wire2202 = {5'd4, 5'd3};
    assign wire2203 = {5'd4, 5'd3};
    assign wire2204 = {5'd4, 5'd3};
    assign wire2205 = {5'd4, 5'd3};
    assign wire2206 = {5'd4, 5'd3};
    assign wire2207 = {5'd4, 5'd3};
    assign wire2208 = {5'd5, 5'd3};
    assign wire2209 = {5'd5, 5'd3};
    assign wire2210 = {5'd5, 5'd3};
    assign wire2211 = {5'd5, 5'd3};
    assign wire2212 = {5'd6, 5'd4};
    assign wire2213 = {5'd9, 5'd7};
    assign wire2214 = {5'd5, 5'd3};
    assign wire2215 = {5'd5, 5'd3};
    assign wire2216 = {5'd6, 5'd4};
    assign wire2217 = {5'd6, 5'd4};
    assign wire2218 = {5'd6, 5'd4};
    assign wire2219 = {5'd6, 5'd4};
    assign wire2220 = {5'd7, 5'd5};
    assign wire2221 = {5'd6, 5'd4};
    assign wire2222 = {5'd6, 5'd4};
    assign wire2223 = {5'd6, 5'd4};
    assign wire2224 = {5'd9, 5'd7};
    assign wire2225 = {5'd9, 5'd7};
    assign wire2226 = {5'd9, 5'd7};
    assign wire2227 = {5'd9, 5'd7};
    assign wire2228 = {5'd10, 5'd8};
    assign wire2229 = {5'd9, 5'd7};
    assign wire2230 = {5'd9, 5'd7};
    assign wire2231 = {5'd9, 5'd7};
    assign wire2232 = {5'd5, 5'd3};
    assign wire2233 = {5'd5, 5'd3};
    assign wire2234 = {5'd5, 5'd3};
    assign wire2235 = {5'd5, 5'd3};
    assign wire2236 = {5'd5, 5'd3};
    assign wire2237 = {5'd5, 5'd3};
    assign wire2238 = {5'd5, 5'd3};
    assign wire2239 = {5'd5, 5'd3};
    assign wire2240 = {5'd7, 5'd3};
    assign wire2241 = {5'd7, 5'd3};
    assign wire2242 = {5'd7, 5'd3};
    assign wire2243 = {5'd7, 5'd3};
    assign wire2244 = {5'd8, 5'd4};
    assign wire2245 = {5'd11, 5'd7};
    assign wire2246 = {5'd7, 5'd3};
    assign wire2247 = {5'd7, 5'd3};
    assign wire2248 = {5'd8, 5'd4};
    assign wire2249 = {5'd8, 5'd4};
    assign wire2250 = {5'd8, 5'd4};
    assign wire2251 = {5'd8, 5'd4};
    assign wire2252 = {5'd9, 5'd5};
    assign wire2253 = {5'd8, 5'd4};
    assign wire2254 = {5'd8, 5'd4};
    assign wire2255 = {5'd8, 5'd4};
    assign wire2256 = {5'd11, 5'd7};
    assign wire2257 = {5'd11, 5'd7};
    assign wire2258 = {5'd11, 5'd7};
    assign wire2259 = {5'd11, 5'd7};
    assign wire2260 = {5'd12, 5'd8};
    assign wire2261 = {5'd11, 5'd7};
    assign wire2262 = {5'd11, 5'd7};
    assign wire2263 = {5'd11, 5'd7};
    assign wire2264 = {5'd7, 5'd3};
    assign wire2265 = {5'd7, 5'd3};
    assign wire2266 = {5'd7, 5'd3};
    assign wire2267 = {5'd7, 5'd3};
    assign wire2268 = {5'd7, 5'd3};
    assign wire2269 = {5'd7, 5'd3};
    assign wire2270 = {5'd7, 5'd3};
    assign wire2271 = {5'd7, 5'd3};
    assign wire2272 = {5'd9, 5'd3};
    assign wire2273 = {5'd9, 5'd3};
    assign wire2274 = {5'd9, 5'd3};
    assign wire2275 = {5'd9, 5'd3};
    assign wire2276 = {5'd10, 5'd4};
    assign wire2277 = {5'd13, 5'd7};
    assign wire2278 = {5'd9, 5'd3};
    assign wire2279 = {5'd9, 5'd3};
    assign wire2280 = {5'd10, 5'd4};
    assign wire2281 = {5'd10, 5'd4};
    assign wire2282 = {5'd10, 5'd4};
    assign wire2283 = {5'd10, 5'd4};
    assign wire2284 = {5'd11, 5'd5};
    assign wire2285 = {5'd10, 5'd4};
    assign wire2286 = {5'd10, 5'd4};
    assign wire2287 = {5'd10, 5'd4};
    assign wire2288 = {5'd13, 5'd7};
    assign wire2289 = {5'd13, 5'd7};
    assign wire2290 = {5'd13, 5'd7};
    assign wire2291 = {5'd13, 5'd7};
    assign wire2292 = {5'd14, 5'd8};
    assign wire2293 = {5'd13, 5'd7};
    assign wire2294 = {5'd13, 5'd7};
    assign wire2295 = {5'd13, 5'd7};
    assign wire2296 = {5'd9, 5'd3};
    assign wire2297 = {5'd9, 5'd3};
    assign wire2298 = {5'd9, 5'd3};
    assign wire2299 = {5'd9, 5'd3};
    assign wire2300 = {5'd9, 5'd3};
    assign wire2301 = {5'd9, 5'd3};
    assign wire2302 = {5'd9, 5'd3};
    assign wire2303 = {5'd9, 5'd3};
    assign wire2304 = {5'd4, 5'd3};
    assign wire2305 = {5'd4, 5'd3};
    assign wire2306 = {5'd4, 5'd3};
    assign wire2307 = {5'd4, 5'd3};
    assign wire2308 = {5'd4, 5'd3};
    assign wire2309 = {5'd4, 5'd3};
    assign wire2310 = {5'd4, 5'd3};
    assign wire2311 = {5'd4, 5'd3};
    assign wire2312 = {5'd4, 5'd3};
    assign wire2313 = {5'd4, 5'd3};
    assign wire2314 = {5'd4, 5'd3};
    assign wire2315 = {5'd4, 5'd3};
    assign wire2316 = {5'd4, 5'd3};
    assign wire2317 = {5'd4, 5'd3};
    assign wire2318 = {5'd4, 5'd3};
    assign wire2319 = {5'd4, 5'd3};
    assign wire2320 = {5'd4, 5'd3};
    assign wire2321 = {5'd4, 5'd3};
    assign wire2322 = {5'd4, 5'd3};
    assign wire2323 = {5'd4, 5'd3};
    assign wire2324 = {5'd4, 5'd3};
    assign wire2325 = {5'd4, 5'd3};
    assign wire2326 = {5'd4, 5'd3};
    assign wire2327 = {5'd4, 5'd3};
    assign wire2328 = {5'd4, 5'd3};
    assign wire2329 = {5'd4, 5'd3};
    assign wire2330 = {5'd4, 5'd3};
    assign wire2331 = {5'd4, 5'd3};
    assign wire2332 = {5'd4, 5'd3};
    assign wire2333 = {5'd4, 5'd3};
    assign wire2334 = {5'd4, 5'd3};
    assign wire2335 = {5'd4, 5'd3};
    assign wire2336 = {5'd5, 5'd3};
    assign wire2337 = {5'd5, 5'd3};
    assign wire2338 = {5'd5, 5'd3};
    assign wire2339 = {5'd5, 5'd3};
    assign wire2340 = {5'd5, 5'd3};
    assign wire2341 = {5'd5, 5'd3};
    assign wire2342 = {5'd5, 5'd3};
    assign wire2343 = {5'd5, 5'd3};
    assign wire2344 = {5'd5, 5'd3};
    assign wire2345 = {5'd5, 5'd3};
    assign wire2346 = {5'd5, 5'd3};
    assign wire2347 = {5'd5, 5'd3};
    assign wire2348 = {5'd5, 5'd3};
    assign wire2349 = {5'd5, 5'd3};
    assign wire2350 = {5'd5, 5'd3};
    assign wire2351 = {5'd5, 5'd3};
    assign wire2352 = {5'd5, 5'd3};
    assign wire2353 = {5'd5, 5'd3};
    assign wire2354 = {5'd5, 5'd3};
    assign wire2355 = {5'd5, 5'd3};
    assign wire2356 = {5'd5, 5'd3};
    assign wire2357 = {5'd5, 5'd3};
    assign wire2358 = {5'd5, 5'd3};
    assign wire2359 = {5'd5, 5'd3};
    assign wire2360 = {5'd5, 5'd3};
    assign wire2361 = {5'd5, 5'd3};
    assign wire2362 = {5'd5, 5'd3};
    assign wire2363 = {5'd5, 5'd3};
    assign wire2364 = {5'd5, 5'd3};
    assign wire2365 = {5'd5, 5'd3};
    assign wire2366 = {5'd5, 5'd3};
    assign wire2367 = {5'd5, 5'd3};
    assign wire2368 = {5'd7, 5'd3};
    assign wire2369 = {5'd7, 5'd3};
    assign wire2370 = {5'd7, 5'd3};
    assign wire2371 = {5'd7, 5'd3};
    assign wire2372 = {5'd7, 5'd3};
    assign wire2373 = {5'd7, 5'd3};
    assign wire2374 = {5'd7, 5'd3};
    assign wire2375 = {5'd7, 5'd3};
    assign wire2376 = {5'd7, 5'd3};
    assign wire2377 = {5'd7, 5'd3};
    assign wire2378 = {5'd7, 5'd3};
    assign wire2379 = {5'd7, 5'd3};
    assign wire2380 = {5'd7, 5'd3};
    assign wire2381 = {5'd7, 5'd3};
    assign wire2382 = {5'd7, 5'd3};
    assign wire2383 = {5'd7, 5'd3};
    assign wire2384 = {5'd7, 5'd3};
    assign wire2385 = {5'd7, 5'd3};
    assign wire2386 = {5'd7, 5'd3};
    assign wire2387 = {5'd7, 5'd3};
    assign wire2388 = {5'd7, 5'd3};
    assign wire2389 = {5'd7, 5'd3};
    assign wire2390 = {5'd7, 5'd3};
    assign wire2391 = {5'd7, 5'd3};
    assign wire2392 = {5'd7, 5'd3};
    assign wire2393 = {5'd7, 5'd3};
    assign wire2394 = {5'd7, 5'd3};
    assign wire2395 = {5'd7, 5'd3};
    assign wire2396 = {5'd7, 5'd3};
    assign wire2397 = {5'd7, 5'd3};
    assign wire2398 = {5'd7, 5'd3};
    assign wire2399 = {5'd7, 5'd3};
    assign wire2400 = {5'd9, 5'd3};
    assign wire2401 = {5'd9, 5'd3};
    assign wire2402 = {5'd9, 5'd3};
    assign wire2403 = {5'd9, 5'd3};
    assign wire2404 = {5'd9, 5'd3};
    assign wire2405 = {5'd9, 5'd3};
    assign wire2406 = {5'd9, 5'd3};
    assign wire2407 = {5'd9, 5'd3};
    assign wire2408 = {5'd9, 5'd3};
    assign wire2409 = {5'd9, 5'd3};
    assign wire2410 = {5'd9, 5'd3};
    assign wire2411 = {5'd9, 5'd3};
    assign wire2412 = {5'd9, 5'd3};
    assign wire2413 = {5'd9, 5'd3};
    assign wire2414 = {5'd9, 5'd3};
    assign wire2415 = {5'd9, 5'd3};
    assign wire2416 = {5'd9, 5'd3};
    assign wire2417 = {5'd9, 5'd3};
    assign wire2418 = {5'd9, 5'd3};
    assign wire2419 = {5'd9, 5'd3};
    assign wire2420 = {5'd9, 5'd3};
    assign wire2421 = {5'd9, 5'd3};
    assign wire2422 = {5'd9, 5'd3};
    assign wire2423 = {5'd9, 5'd3};
    assign wire2424 = {5'd9, 5'd3};
    assign wire2425 = {5'd9, 5'd3};
    assign wire2426 = {5'd9, 5'd3};
    assign wire2427 = {5'd9, 5'd3};
    assign wire2428 = {5'd9, 5'd3};
    assign wire2429 = {5'd9, 5'd3};
    assign wire2430 = {5'd9, 5'd3};
    assign wire2431 = {5'd9, 5'd3};
    assign wire2432 = {5'd5, 5'd4};
    assign wire2433 = {5'd5, 5'd4};
    assign wire2434 = {5'd5, 5'd4};
    assign wire2435 = {5'd5, 5'd4};
    assign wire2436 = {5'd6, 5'd5};
    assign wire2437 = {5'd9, 5'd8};
    assign wire2438 = {5'd5, 5'd4};
    assign wire2439 = {5'd5, 5'd4};
    assign wire2440 = {5'd6, 5'd5};
    assign wire2441 = {5'd6, 5'd5};
    assign wire2442 = {5'd6, 5'd5};
    assign wire2443 = {5'd6, 5'd5};
    assign wire2444 = {5'd7, 5'd6};
    assign wire2445 = {5'd6, 5'd5};
    assign wire2446 = {5'd6, 5'd5};
    assign wire2447 = {5'd6, 5'd5};
    assign wire2448 = {5'd9, 5'd8};
    assign wire2449 = {5'd9, 5'd8};
    assign wire2450 = {5'd9, 5'd8};
    assign wire2451 = {5'd9, 5'd8};
    assign wire2452 = {5'd10, 5'd9};
    assign wire2453 = {5'd9, 5'd8};
    assign wire2454 = {5'd9, 5'd8};
    assign wire2455 = {5'd9, 5'd8};
    assign wire2456 = {5'd5, 5'd4};
    assign wire2457 = {5'd5, 5'd4};
    assign wire2458 = {5'd5, 5'd4};
    assign wire2459 = {5'd5, 5'd4};
    assign wire2460 = {5'd5, 5'd4};
    assign wire2461 = {5'd5, 5'd4};
    assign wire2462 = {5'd5, 5'd4};
    assign wire2463 = {5'd5, 5'd4};
    assign wire2464 = {5'd6, 5'd4};
    assign wire2465 = {5'd6, 5'd4};
    assign wire2466 = {5'd6, 5'd4};
    assign wire2467 = {5'd6, 5'd4};
    assign wire2468 = {5'd7, 5'd5};
    assign wire2469 = {5'd10, 5'd8};
    assign wire2470 = {5'd6, 5'd4};
    assign wire2471 = {5'd6, 5'd4};
    assign wire2472 = {5'd7, 5'd5};
    assign wire2473 = {5'd7, 5'd5};
    assign wire2474 = {5'd7, 5'd5};
    assign wire2475 = {5'd7, 5'd5};
    assign wire2476 = {5'd8, 5'd6};
    assign wire2477 = {5'd7, 5'd5};
    assign wire2478 = {5'd7, 5'd5};
    assign wire2479 = {5'd7, 5'd5};
    assign wire2480 = {5'd10, 5'd8};
    assign wire2481 = {5'd10, 5'd8};
    assign wire2482 = {5'd10, 5'd8};
    assign wire2483 = {5'd10, 5'd8};
    assign wire2484 = {5'd11, 5'd9};
    assign wire2485 = {5'd10, 5'd8};
    assign wire2486 = {5'd10, 5'd8};
    assign wire2487 = {5'd10, 5'd8};
    assign wire2488 = {5'd6, 5'd4};
    assign wire2489 = {5'd6, 5'd4};
    assign wire2490 = {5'd6, 5'd4};
    assign wire2491 = {5'd6, 5'd4};
    assign wire2492 = {5'd6, 5'd4};
    assign wire2493 = {5'd6, 5'd4};
    assign wire2494 = {5'd6, 5'd4};
    assign wire2495 = {5'd6, 5'd4};
    assign wire2496 = {5'd8, 5'd4};
    assign wire2497 = {5'd8, 5'd4};
    assign wire2498 = {5'd8, 5'd4};
    assign wire2499 = {5'd8, 5'd4};
    assign wire2500 = {5'd9, 5'd5};
    assign wire2501 = {5'd12, 5'd8};
    assign wire2502 = {5'd8, 5'd4};
    assign wire2503 = {5'd8, 5'd4};
    assign wire2504 = {5'd9, 5'd5};
    assign wire2505 = {5'd9, 5'd5};
    assign wire2506 = {5'd9, 5'd5};
    assign wire2507 = {5'd9, 5'd5};
    assign wire2508 = {5'd10, 5'd6};
    assign wire2509 = {5'd9, 5'd5};
    assign wire2510 = {5'd9, 5'd5};
    assign wire2511 = {5'd9, 5'd5};
    assign wire2512 = {5'd12, 5'd8};
    assign wire2513 = {5'd12, 5'd8};
    assign wire2514 = {5'd12, 5'd8};
    assign wire2515 = {5'd12, 5'd8};
    assign wire2516 = {5'd13, 5'd9};
    assign wire2517 = {5'd12, 5'd8};
    assign wire2518 = {5'd12, 5'd8};
    assign wire2519 = {5'd12, 5'd8};
    assign wire2520 = {5'd8, 5'd4};
    assign wire2521 = {5'd8, 5'd4};
    assign wire2522 = {5'd8, 5'd4};
    assign wire2523 = {5'd8, 5'd4};
    assign wire2524 = {5'd8, 5'd4};
    assign wire2525 = {5'd8, 5'd4};
    assign wire2526 = {5'd8, 5'd4};
    assign wire2527 = {5'd8, 5'd4};
    assign wire2528 = {5'd10, 5'd4};
    assign wire2529 = {5'd10, 5'd4};
    assign wire2530 = {5'd10, 5'd4};
    assign wire2531 = {5'd10, 5'd4};
    assign wire2532 = {5'd11, 5'd5};
    assign wire2533 = {5'd14, 5'd8};
    assign wire2534 = {5'd10, 5'd4};
    assign wire2535 = {5'd10, 5'd4};
    assign wire2536 = {5'd11, 5'd5};
    assign wire2537 = {5'd11, 5'd5};
    assign wire2538 = {5'd11, 5'd5};
    assign wire2539 = {5'd11, 5'd5};
    assign wire2540 = {5'd12, 5'd6};
    assign wire2541 = {5'd11, 5'd5};
    assign wire2542 = {5'd11, 5'd5};
    assign wire2543 = {5'd11, 5'd5};
    assign wire2544 = {5'd14, 5'd8};
    assign wire2545 = {5'd14, 5'd8};
    assign wire2546 = {5'd14, 5'd8};
    assign wire2547 = {5'd14, 5'd8};
    assign wire2548 = {5'd15, 5'd9};
    assign wire2549 = {5'd14, 5'd8};
    assign wire2550 = {5'd14, 5'd8};
    assign wire2551 = {5'd14, 5'd8};
    assign wire2552 = {5'd10, 5'd4};
    assign wire2553 = {5'd10, 5'd4};
    assign wire2554 = {5'd10, 5'd4};
    assign wire2555 = {5'd10, 5'd4};
    assign wire2556 = {5'd10, 5'd4};
    assign wire2557 = {5'd10, 5'd4};
    assign wire2558 = {5'd10, 5'd4};
    assign wire2559 = {5'd10, 5'd4};
    assign wire2560 = {5'd4, 5'd3};
    assign wire2561 = {5'd4, 5'd3};
    assign wire2562 = {5'd4, 5'd3};
    assign wire2563 = {5'd4, 5'd3};
    assign wire2564 = {5'd4, 5'd3};
    assign wire2565 = {5'd4, 5'd3};
    assign wire2566 = {5'd4, 5'd3};
    assign wire2567 = {5'd4, 5'd3};
    assign wire2568 = {5'd4, 5'd3};
    assign wire2569 = {5'd4, 5'd3};
    assign wire2570 = {5'd4, 5'd3};
    assign wire2571 = {5'd4, 5'd3};
    assign wire2572 = {5'd4, 5'd3};
    assign wire2573 = {5'd4, 5'd3};
    assign wire2574 = {5'd4, 5'd3};
    assign wire2575 = {5'd4, 5'd3};
    assign wire2576 = {5'd4, 5'd3};
    assign wire2577 = {5'd4, 5'd3};
    assign wire2578 = {5'd4, 5'd3};
    assign wire2579 = {5'd4, 5'd3};
    assign wire2580 = {5'd4, 5'd3};
    assign wire2581 = {5'd4, 5'd3};
    assign wire2582 = {5'd4, 5'd3};
    assign wire2583 = {5'd4, 5'd3};
    assign wire2584 = {5'd4, 5'd3};
    assign wire2585 = {5'd4, 5'd3};
    assign wire2586 = {5'd4, 5'd3};
    assign wire2587 = {5'd4, 5'd3};
    assign wire2588 = {5'd4, 5'd3};
    assign wire2589 = {5'd4, 5'd3};
    assign wire2590 = {5'd4, 5'd3};
    assign wire2591 = {5'd4, 5'd3};
    assign wire2592 = {5'd5, 5'd3};
    assign wire2593 = {5'd5, 5'd3};
    assign wire2594 = {5'd5, 5'd3};
    assign wire2595 = {5'd5, 5'd3};
    assign wire2596 = {5'd5, 5'd3};
    assign wire2597 = {5'd5, 5'd3};
    assign wire2598 = {5'd5, 5'd3};
    assign wire2599 = {5'd5, 5'd3};
    assign wire2600 = {5'd5, 5'd3};
    assign wire2601 = {5'd5, 5'd3};
    assign wire2602 = {5'd5, 5'd3};
    assign wire2603 = {5'd5, 5'd3};
    assign wire2604 = {5'd5, 5'd3};
    assign wire2605 = {5'd5, 5'd3};
    assign wire2606 = {5'd5, 5'd3};
    assign wire2607 = {5'd5, 5'd3};
    assign wire2608 = {5'd5, 5'd3};
    assign wire2609 = {5'd5, 5'd3};
    assign wire2610 = {5'd5, 5'd3};
    assign wire2611 = {5'd5, 5'd3};
    assign wire2612 = {5'd5, 5'd3};
    assign wire2613 = {5'd5, 5'd3};
    assign wire2614 = {5'd5, 5'd3};
    assign wire2615 = {5'd5, 5'd3};
    assign wire2616 = {5'd5, 5'd3};
    assign wire2617 = {5'd5, 5'd3};
    assign wire2618 = {5'd5, 5'd3};
    assign wire2619 = {5'd5, 5'd3};
    assign wire2620 = {5'd5, 5'd3};
    assign wire2621 = {5'd5, 5'd3};
    assign wire2622 = {5'd5, 5'd3};
    assign wire2623 = {5'd5, 5'd3};
    assign wire2624 = {5'd7, 5'd3};
    assign wire2625 = {5'd7, 5'd3};
    assign wire2626 = {5'd7, 5'd3};
    assign wire2627 = {5'd7, 5'd3};
    assign wire2628 = {5'd7, 5'd3};
    assign wire2629 = {5'd7, 5'd3};
    assign wire2630 = {5'd7, 5'd3};
    assign wire2631 = {5'd7, 5'd3};
    assign wire2632 = {5'd7, 5'd3};
    assign wire2633 = {5'd7, 5'd3};
    assign wire2634 = {5'd7, 5'd3};
    assign wire2635 = {5'd7, 5'd3};
    assign wire2636 = {5'd7, 5'd3};
    assign wire2637 = {5'd7, 5'd3};
    assign wire2638 = {5'd7, 5'd3};
    assign wire2639 = {5'd7, 5'd3};
    assign wire2640 = {5'd7, 5'd3};
    assign wire2641 = {5'd7, 5'd3};
    assign wire2642 = {5'd7, 5'd3};
    assign wire2643 = {5'd7, 5'd3};
    assign wire2644 = {5'd7, 5'd3};
    assign wire2645 = {5'd7, 5'd3};
    assign wire2646 = {5'd7, 5'd3};
    assign wire2647 = {5'd7, 5'd3};
    assign wire2648 = {5'd7, 5'd3};
    assign wire2649 = {5'd7, 5'd3};
    assign wire2650 = {5'd7, 5'd3};
    assign wire2651 = {5'd7, 5'd3};
    assign wire2652 = {5'd7, 5'd3};
    assign wire2653 = {5'd7, 5'd3};
    assign wire2654 = {5'd7, 5'd3};
    assign wire2655 = {5'd7, 5'd3};
    assign wire2656 = {5'd9, 5'd3};
    assign wire2657 = {5'd9, 5'd3};
    assign wire2658 = {5'd9, 5'd3};
    assign wire2659 = {5'd9, 5'd3};
    assign wire2660 = {5'd9, 5'd3};
    assign wire2661 = {5'd9, 5'd3};
    assign wire2662 = {5'd9, 5'd3};
    assign wire2663 = {5'd9, 5'd3};
    assign wire2664 = {5'd9, 5'd3};
    assign wire2665 = {5'd9, 5'd3};
    assign wire2666 = {5'd9, 5'd3};
    assign wire2667 = {5'd9, 5'd3};
    assign wire2668 = {5'd9, 5'd3};
    assign wire2669 = {5'd9, 5'd3};
    assign wire2670 = {5'd9, 5'd3};
    assign wire2671 = {5'd9, 5'd3};
    assign wire2672 = {5'd9, 5'd3};
    assign wire2673 = {5'd9, 5'd3};
    assign wire2674 = {5'd9, 5'd3};
    assign wire2675 = {5'd9, 5'd3};
    assign wire2676 = {5'd9, 5'd3};
    assign wire2677 = {5'd9, 5'd3};
    assign wire2678 = {5'd9, 5'd3};
    assign wire2679 = {5'd9, 5'd3};
    assign wire2680 = {5'd9, 5'd3};
    assign wire2681 = {5'd9, 5'd3};
    assign wire2682 = {5'd9, 5'd3};
    assign wire2683 = {5'd9, 5'd3};
    assign wire2684 = {5'd9, 5'd3};
    assign wire2685 = {5'd9, 5'd3};
    assign wire2686 = {5'd9, 5'd3};
    assign wire2687 = {5'd9, 5'd3};
    assign wire2688 = {5'd5, 5'd4};
    assign wire2689 = {5'd5, 5'd4};
    assign wire2690 = {5'd5, 5'd4};
    assign wire2691 = {5'd5, 5'd4};
    assign wire2692 = {5'd5, 5'd4};
    assign wire2693 = {5'd7, 5'd6};
    assign wire2694 = {5'd5, 5'd4};
    assign wire2695 = {5'd5, 5'd4};
    assign wire2696 = {5'd6, 5'd5};
    assign wire2697 = {5'd6, 5'd5};
    assign wire2698 = {5'd6, 5'd5};
    assign wire2699 = {5'd6, 5'd5};
    assign wire2700 = {5'd6, 5'd5};
    assign wire2701 = {5'd6, 5'd5};
    assign wire2702 = {5'd6, 5'd5};
    assign wire2703 = {5'd6, 5'd5};
    assign wire2704 = {5'd7, 5'd6};
    assign wire2705 = {5'd7, 5'd6};
    assign wire2706 = {5'd7, 5'd6};
    assign wire2707 = {5'd7, 5'd6};
    assign wire2708 = {5'd7, 5'd6};
    assign wire2709 = {5'd7, 5'd6};
    assign wire2710 = {5'd7, 5'd6};
    assign wire2711 = {5'd7, 5'd6};
    assign wire2712 = {5'd5, 5'd4};
    assign wire2713 = {5'd5, 5'd4};
    assign wire2714 = {5'd5, 5'd4};
    assign wire2715 = {5'd5, 5'd4};
    assign wire2716 = {5'd5, 5'd4};
    assign wire2717 = {5'd5, 5'd4};
    assign wire2718 = {5'd5, 5'd4};
    assign wire2719 = {5'd5, 5'd4};
    assign wire2720 = {5'd6, 5'd4};
    assign wire2721 = {5'd6, 5'd4};
    assign wire2722 = {5'd6, 5'd4};
    assign wire2723 = {5'd6, 5'd4};
    assign wire2724 = {5'd6, 5'd4};
    assign wire2725 = {5'd8, 5'd6};
    assign wire2726 = {5'd6, 5'd4};
    assign wire2727 = {5'd6, 5'd4};
    assign wire2728 = {5'd7, 5'd5};
    assign wire2729 = {5'd7, 5'd5};
    assign wire2730 = {5'd7, 5'd5};
    assign wire2731 = {5'd7, 5'd5};
    assign wire2732 = {5'd7, 5'd5};
    assign wire2733 = {5'd7, 5'd5};
    assign wire2734 = {5'd7, 5'd5};
    assign wire2735 = {5'd7, 5'd5};
    assign wire2736 = {5'd8, 5'd6};
    assign wire2737 = {5'd8, 5'd6};
    assign wire2738 = {5'd8, 5'd6};
    assign wire2739 = {5'd8, 5'd6};
    assign wire2740 = {5'd8, 5'd6};
    assign wire2741 = {5'd8, 5'd6};
    assign wire2742 = {5'd8, 5'd6};
    assign wire2743 = {5'd8, 5'd6};
    assign wire2744 = {5'd6, 5'd4};
    assign wire2745 = {5'd6, 5'd4};
    assign wire2746 = {5'd6, 5'd4};
    assign wire2747 = {5'd6, 5'd4};
    assign wire2748 = {5'd6, 5'd4};
    assign wire2749 = {5'd6, 5'd4};
    assign wire2750 = {5'd6, 5'd4};
    assign wire2751 = {5'd6, 5'd4};
    assign wire2752 = {5'd8, 5'd4};
    assign wire2753 = {5'd8, 5'd4};
    assign wire2754 = {5'd8, 5'd4};
    assign wire2755 = {5'd8, 5'd4};
    assign wire2756 = {5'd8, 5'd4};
    assign wire2757 = {5'd10, 5'd6};
    assign wire2758 = {5'd8, 5'd4};
    assign wire2759 = {5'd8, 5'd4};
    assign wire2760 = {5'd9, 5'd5};
    assign wire2761 = {5'd9, 5'd5};
    assign wire2762 = {5'd9, 5'd5};
    assign wire2763 = {5'd9, 5'd5};
    assign wire2764 = {5'd9, 5'd5};
    assign wire2765 = {5'd9, 5'd5};
    assign wire2766 = {5'd9, 5'd5};
    assign wire2767 = {5'd9, 5'd5};
    assign wire2768 = {5'd10, 5'd6};
    assign wire2769 = {5'd10, 5'd6};
    assign wire2770 = {5'd10, 5'd6};
    assign wire2771 = {5'd10, 5'd6};
    assign wire2772 = {5'd10, 5'd6};
    assign wire2773 = {5'd10, 5'd6};
    assign wire2774 = {5'd10, 5'd6};
    assign wire2775 = {5'd10, 5'd6};
    assign wire2776 = {5'd8, 5'd4};
    assign wire2777 = {5'd8, 5'd4};
    assign wire2778 = {5'd8, 5'd4};
    assign wire2779 = {5'd8, 5'd4};
    assign wire2780 = {5'd8, 5'd4};
    assign wire2781 = {5'd8, 5'd4};
    assign wire2782 = {5'd8, 5'd4};
    assign wire2783 = {5'd8, 5'd4};
    assign wire2784 = {5'd10, 5'd4};
    assign wire2785 = {5'd10, 5'd4};
    assign wire2786 = {5'd10, 5'd4};
    assign wire2787 = {5'd10, 5'd4};
    assign wire2788 = {5'd10, 5'd4};
    assign wire2789 = {5'd12, 5'd6};
    assign wire2790 = {5'd10, 5'd4};
    assign wire2791 = {5'd10, 5'd4};
    assign wire2792 = {5'd11, 5'd5};
    assign wire2793 = {5'd11, 5'd5};
    assign wire2794 = {5'd11, 5'd5};
    assign wire2795 = {5'd11, 5'd5};
    assign wire2796 = {5'd11, 5'd5};
    assign wire2797 = {5'd11, 5'd5};
    assign wire2798 = {5'd11, 5'd5};
    assign wire2799 = {5'd11, 5'd5};
    assign wire2800 = {5'd12, 5'd6};
    assign wire2801 = {5'd12, 5'd6};
    assign wire2802 = {5'd12, 5'd6};
    assign wire2803 = {5'd12, 5'd6};
    assign wire2804 = {5'd12, 5'd6};
    assign wire2805 = {5'd12, 5'd6};
    assign wire2806 = {5'd12, 5'd6};
    assign wire2807 = {5'd12, 5'd6};
    assign wire2808 = {5'd10, 5'd4};
    assign wire2809 = {5'd10, 5'd4};
    assign wire2810 = {5'd10, 5'd4};
    assign wire2811 = {5'd10, 5'd4};
    assign wire2812 = {5'd10, 5'd4};
    assign wire2813 = {5'd10, 5'd4};
    assign wire2814 = {5'd10, 5'd4};
    assign wire2815 = {5'd10, 5'd4};
    assign wire2816 = {5'd5, 5'd4};
    assign wire2817 = {5'd5, 5'd4};
    assign wire2818 = {5'd5, 5'd4};
    assign wire2819 = {5'd5, 5'd4};
    assign wire2820 = {5'd5, 5'd4};
    assign wire2821 = {5'd5, 5'd4};
    assign wire2822 = {5'd5, 5'd4};
    assign wire2823 = {5'd5, 5'd4};
    assign wire2824 = {5'd5, 5'd4};
    assign wire2825 = {5'd5, 5'd4};
    assign wire2826 = {5'd5, 5'd4};
    assign wire2827 = {5'd5, 5'd4};
    assign wire2828 = {5'd5, 5'd4};
    assign wire2829 = {5'd5, 5'd4};
    assign wire2830 = {5'd5, 5'd4};
    assign wire2831 = {5'd5, 5'd4};
    assign wire2832 = {5'd5, 5'd4};
    assign wire2833 = {5'd5, 5'd4};
    assign wire2834 = {5'd5, 5'd4};
    assign wire2835 = {5'd5, 5'd4};
    assign wire2836 = {5'd5, 5'd4};
    assign wire2837 = {5'd5, 5'd4};
    assign wire2838 = {5'd5, 5'd4};
    assign wire2839 = {5'd5, 5'd4};
    assign wire2840 = {5'd5, 5'd4};
    assign wire2841 = {5'd5, 5'd4};
    assign wire2842 = {5'd5, 5'd4};
    assign wire2843 = {5'd5, 5'd4};
    assign wire2844 = {5'd5, 5'd4};
    assign wire2845 = {5'd5, 5'd4};
    assign wire2846 = {5'd5, 5'd4};
    assign wire2847 = {5'd5, 5'd4};
    assign wire2848 = {5'd6, 5'd4};
    assign wire2849 = {5'd6, 5'd4};
    assign wire2850 = {5'd6, 5'd4};
    assign wire2851 = {5'd6, 5'd4};
    assign wire2852 = {5'd6, 5'd4};
    assign wire2853 = {5'd6, 5'd4};
    assign wire2854 = {5'd6, 5'd4};
    assign wire2855 = {5'd6, 5'd4};
    assign wire2856 = {5'd6, 5'd4};
    assign wire2857 = {5'd6, 5'd4};
    assign wire2858 = {5'd6, 5'd4};
    assign wire2859 = {5'd6, 5'd4};
    assign wire2860 = {5'd6, 5'd4};
    assign wire2861 = {5'd6, 5'd4};
    assign wire2862 = {5'd6, 5'd4};
    assign wire2863 = {5'd6, 5'd4};
    assign wire2864 = {5'd6, 5'd4};
    assign wire2865 = {5'd6, 5'd4};
    assign wire2866 = {5'd6, 5'd4};
    assign wire2867 = {5'd6, 5'd4};
    assign wire2868 = {5'd6, 5'd4};
    assign wire2869 = {5'd6, 5'd4};
    assign wire2870 = {5'd6, 5'd4};
    assign wire2871 = {5'd6, 5'd4};
    assign wire2872 = {5'd6, 5'd4};
    assign wire2873 = {5'd6, 5'd4};
    assign wire2874 = {5'd6, 5'd4};
    assign wire2875 = {5'd6, 5'd4};
    assign wire2876 = {5'd6, 5'd4};
    assign wire2877 = {5'd6, 5'd4};
    assign wire2878 = {5'd6, 5'd4};
    assign wire2879 = {5'd6, 5'd4};
    assign wire2880 = {5'd8, 5'd4};
    assign wire2881 = {5'd8, 5'd4};
    assign wire2882 = {5'd8, 5'd4};
    assign wire2883 = {5'd8, 5'd4};
    assign wire2884 = {5'd8, 5'd4};
    assign wire2885 = {5'd8, 5'd4};
    assign wire2886 = {5'd8, 5'd4};
    assign wire2887 = {5'd8, 5'd4};
    assign wire2888 = {5'd8, 5'd4};
    assign wire2889 = {5'd8, 5'd4};
    assign wire2890 = {5'd8, 5'd4};
    assign wire2891 = {5'd8, 5'd4};
    assign wire2892 = {5'd8, 5'd4};
    assign wire2893 = {5'd8, 5'd4};
    assign wire2894 = {5'd8, 5'd4};
    assign wire2895 = {5'd8, 5'd4};
    assign wire2896 = {5'd8, 5'd4};
    assign wire2897 = {5'd8, 5'd4};
    assign wire2898 = {5'd8, 5'd4};
    assign wire2899 = {5'd8, 5'd4};
    assign wire2900 = {5'd8, 5'd4};
    assign wire2901 = {5'd8, 5'd4};
    assign wire2902 = {5'd8, 5'd4};
    assign wire2903 = {5'd8, 5'd4};
    assign wire2904 = {5'd8, 5'd4};
    assign wire2905 = {5'd8, 5'd4};
    assign wire2906 = {5'd8, 5'd4};
    assign wire2907 = {5'd8, 5'd4};
    assign wire2908 = {5'd8, 5'd4};
    assign wire2909 = {5'd8, 5'd4};
    assign wire2910 = {5'd8, 5'd4};
    assign wire2911 = {5'd8, 5'd4};
    assign wire2912 = {5'd10, 5'd4};
    assign wire2913 = {5'd10, 5'd4};
    assign wire2914 = {5'd10, 5'd4};
    assign wire2915 = {5'd10, 5'd4};
    assign wire2916 = {5'd10, 5'd4};
    assign wire2917 = {5'd10, 5'd4};
    assign wire2918 = {5'd10, 5'd4};
    assign wire2919 = {5'd10, 5'd4};
    assign wire2920 = {5'd10, 5'd4};
    assign wire2921 = {5'd10, 5'd4};
    assign wire2922 = {5'd10, 5'd4};
    assign wire2923 = {5'd10, 5'd4};
    assign wire2924 = {5'd10, 5'd4};
    assign wire2925 = {5'd10, 5'd4};
    assign wire2926 = {5'd10, 5'd4};
    assign wire2927 = {5'd10, 5'd4};
    assign wire2928 = {5'd10, 5'd4};
    assign wire2929 = {5'd10, 5'd4};
    assign wire2930 = {5'd10, 5'd4};
    assign wire2931 = {5'd10, 5'd4};
    assign wire2932 = {5'd10, 5'd4};
    assign wire2933 = {5'd10, 5'd4};
    assign wire2934 = {5'd10, 5'd4};
    assign wire2935 = {5'd10, 5'd4};
    assign wire2936 = {5'd10, 5'd4};
    assign wire2937 = {5'd10, 5'd4};
    assign wire2938 = {5'd10, 5'd4};
    assign wire2939 = {5'd10, 5'd4};
    assign wire2940 = {5'd10, 5'd4};
    assign wire2941 = {5'd10, 5'd4};
    assign wire2942 = {5'd10, 5'd4};
    assign wire2943 = {5'd10, 5'd4};
    assign wire2944 = {5'd6, 5'd5};
    assign wire2945 = {5'd6, 5'd5};
    assign wire2946 = {5'd6, 5'd5};
    assign wire2947 = {5'd6, 5'd5};
    assign wire2948 = {5'd6, 5'd5};
    assign wire2949 = {5'd8, 5'd7};
    assign wire2950 = {5'd6, 5'd5};
    assign wire2951 = {5'd6, 5'd5};
    assign wire2952 = {5'd7, 5'd6};
    assign wire2953 = {5'd7, 5'd6};
    assign wire2954 = {5'd7, 5'd6};
    assign wire2955 = {5'd7, 5'd6};
    assign wire2956 = {5'd7, 5'd6};
    assign wire2957 = {5'd7, 5'd6};
    assign wire2958 = {5'd7, 5'd6};
    assign wire2959 = {5'd7, 5'd6};
    assign wire2960 = {5'd8, 5'd7};
    assign wire2961 = {5'd8, 5'd7};
    assign wire2962 = {5'd8, 5'd7};
    assign wire2963 = {5'd8, 5'd7};
    assign wire2964 = {5'd8, 5'd7};
    assign wire2965 = {5'd8, 5'd7};
    assign wire2966 = {5'd8, 5'd7};
    assign wire2967 = {5'd8, 5'd7};
    assign wire2968 = {5'd6, 5'd5};
    assign wire2969 = {5'd6, 5'd5};
    assign wire2970 = {5'd6, 5'd5};
    assign wire2971 = {5'd6, 5'd5};
    assign wire2972 = {5'd6, 5'd5};
    assign wire2973 = {5'd6, 5'd5};
    assign wire2974 = {5'd6, 5'd5};
    assign wire2975 = {5'd6, 5'd5};
    assign wire2976 = {5'd7, 5'd5};
    assign wire2977 = {5'd7, 5'd5};
    assign wire2978 = {5'd7, 5'd5};
    assign wire2979 = {5'd7, 5'd5};
    assign wire2980 = {5'd7, 5'd5};
    assign wire2981 = {5'd9, 5'd7};
    assign wire2982 = {5'd7, 5'd5};
    assign wire2983 = {5'd7, 5'd5};
    assign wire2984 = {5'd8, 5'd6};
    assign wire2985 = {5'd8, 5'd6};
    assign wire2986 = {5'd8, 5'd6};
    assign wire2987 = {5'd8, 5'd6};
    assign wire2988 = {5'd8, 5'd6};
    assign wire2989 = {5'd8, 5'd6};
    assign wire2990 = {5'd8, 5'd6};
    assign wire2991 = {5'd8, 5'd6};
    assign wire2992 = {5'd9, 5'd7};
    assign wire2993 = {5'd9, 5'd7};
    assign wire2994 = {5'd9, 5'd7};
    assign wire2995 = {5'd9, 5'd7};
    assign wire2996 = {5'd9, 5'd7};
    assign wire2997 = {5'd9, 5'd7};
    assign wire2998 = {5'd9, 5'd7};
    assign wire2999 = {5'd9, 5'd7};
    assign wire3000 = {5'd7, 5'd5};
    assign wire3001 = {5'd7, 5'd5};
    assign wire3002 = {5'd7, 5'd5};
    assign wire3003 = {5'd7, 5'd5};
    assign wire3004 = {5'd7, 5'd5};
    assign wire3005 = {5'd7, 5'd5};
    assign wire3006 = {5'd7, 5'd5};
    assign wire3007 = {5'd7, 5'd5};
    assign wire3008 = {5'd9, 5'd5};
    assign wire3009 = {5'd9, 5'd5};
    assign wire3010 = {5'd9, 5'd5};
    assign wire3011 = {5'd9, 5'd5};
    assign wire3012 = {5'd9, 5'd5};
    assign wire3013 = {5'd11, 5'd7};
    assign wire3014 = {5'd9, 5'd5};
    assign wire3015 = {5'd9, 5'd5};
    assign wire3016 = {5'd10, 5'd6};
    assign wire3017 = {5'd10, 5'd6};
    assign wire3018 = {5'd10, 5'd6};
    assign wire3019 = {5'd10, 5'd6};
    assign wire3020 = {5'd10, 5'd6};
    assign wire3021 = {5'd10, 5'd6};
    assign wire3022 = {5'd10, 5'd6};
    assign wire3023 = {5'd10, 5'd6};
    assign wire3024 = {5'd11, 5'd7};
    assign wire3025 = {5'd11, 5'd7};
    assign wire3026 = {5'd11, 5'd7};
    assign wire3027 = {5'd11, 5'd7};
    assign wire3028 = {5'd11, 5'd7};
    assign wire3029 = {5'd11, 5'd7};
    assign wire3030 = {5'd11, 5'd7};
    assign wire3031 = {5'd11, 5'd7};
    assign wire3032 = {5'd9, 5'd5};
    assign wire3033 = {5'd9, 5'd5};
    assign wire3034 = {5'd9, 5'd5};
    assign wire3035 = {5'd9, 5'd5};
    assign wire3036 = {5'd9, 5'd5};
    assign wire3037 = {5'd9, 5'd5};
    assign wire3038 = {5'd9, 5'd5};
    assign wire3039 = {5'd9, 5'd5};
    assign wire3040 = {5'd11, 5'd5};
    assign wire3041 = {5'd11, 5'd5};
    assign wire3042 = {5'd11, 5'd5};
    assign wire3043 = {5'd11, 5'd5};
    assign wire3044 = {5'd11, 5'd5};
    assign wire3045 = {5'd13, 5'd7};
    assign wire3046 = {5'd11, 5'd5};
    assign wire3047 = {5'd11, 5'd5};
    assign wire3048 = {5'd12, 5'd6};
    assign wire3049 = {5'd12, 5'd6};
    assign wire3050 = {5'd12, 5'd6};
    assign wire3051 = {5'd12, 5'd6};
    assign wire3052 = {5'd12, 5'd6};
    assign wire3053 = {5'd12, 5'd6};
    assign wire3054 = {5'd12, 5'd6};
    assign wire3055 = {5'd12, 5'd6};
    assign wire3056 = {5'd13, 5'd7};
    assign wire3057 = {5'd13, 5'd7};
    assign wire3058 = {5'd13, 5'd7};
    assign wire3059 = {5'd13, 5'd7};
    assign wire3060 = {5'd13, 5'd7};
    assign wire3061 = {5'd13, 5'd7};
    assign wire3062 = {5'd13, 5'd7};
    assign wire3063 = {5'd13, 5'd7};
    assign wire3064 = {5'd11, 5'd5};
    assign wire3065 = {5'd11, 5'd5};
    assign wire3066 = {5'd11, 5'd5};
    assign wire3067 = {5'd11, 5'd5};
    assign wire3068 = {5'd11, 5'd5};
    assign wire3069 = {5'd11, 5'd5};
    assign wire3070 = {5'd11, 5'd5};
    assign wire3071 = {5'd11, 5'd5};
    assign wire3072 = {5'd4, 5'd3};
    assign wire3073 = {5'd4, 5'd3};
    assign wire3074 = {5'd4, 5'd3};
    assign wire3075 = {5'd4, 5'd3};
    assign wire3076 = {5'd4, 5'd3};
    assign wire3077 = {5'd4, 5'd3};
    assign wire3078 = {5'd4, 5'd3};
    assign wire3079 = {5'd4, 5'd3};
    assign wire3080 = {5'd4, 5'd3};
    assign wire3081 = {5'd4, 5'd3};
    assign wire3082 = {5'd4, 5'd3};
    assign wire3083 = {5'd4, 5'd3};
    assign wire3084 = {5'd4, 5'd3};
    assign wire3085 = {5'd4, 5'd3};
    assign wire3086 = {5'd4, 5'd3};
    assign wire3087 = {5'd4, 5'd3};
    assign wire3088 = {5'd4, 5'd3};
    assign wire3089 = {5'd4, 5'd3};
    assign wire3090 = {5'd4, 5'd3};
    assign wire3091 = {5'd4, 5'd3};
    assign wire3092 = {5'd4, 5'd3};
    assign wire3093 = {5'd4, 5'd3};
    assign wire3094 = {5'd4, 5'd3};
    assign wire3095 = {5'd4, 5'd3};
    assign wire3096 = {5'd4, 5'd3};
    assign wire3097 = {5'd4, 5'd3};
    assign wire3098 = {5'd4, 5'd3};
    assign wire3099 = {5'd4, 5'd3};
    assign wire3100 = {5'd4, 5'd3};
    assign wire3101 = {5'd4, 5'd3};
    assign wire3102 = {5'd4, 5'd3};
    assign wire3103 = {5'd4, 5'd3};
    assign wire3104 = {5'd5, 5'd3};
    assign wire3105 = {5'd5, 5'd3};
    assign wire3106 = {5'd5, 5'd3};
    assign wire3107 = {5'd5, 5'd3};
    assign wire3108 = {5'd5, 5'd3};
    assign wire3109 = {5'd5, 5'd3};
    assign wire3110 = {5'd5, 5'd3};
    assign wire3111 = {5'd5, 5'd3};
    assign wire3112 = {5'd5, 5'd3};
    assign wire3113 = {5'd5, 5'd3};
    assign wire3114 = {5'd5, 5'd3};
    assign wire3115 = {5'd5, 5'd3};
    assign wire3116 = {5'd5, 5'd3};
    assign wire3117 = {5'd5, 5'd3};
    assign wire3118 = {5'd5, 5'd3};
    assign wire3119 = {5'd5, 5'd3};
    assign wire3120 = {5'd5, 5'd3};
    assign wire3121 = {5'd5, 5'd3};
    assign wire3122 = {5'd5, 5'd3};
    assign wire3123 = {5'd5, 5'd3};
    assign wire3124 = {5'd5, 5'd3};
    assign wire3125 = {5'd5, 5'd3};
    assign wire3126 = {5'd5, 5'd3};
    assign wire3127 = {5'd5, 5'd3};
    assign wire3128 = {5'd5, 5'd3};
    assign wire3129 = {5'd5, 5'd3};
    assign wire3130 = {5'd5, 5'd3};
    assign wire3131 = {5'd5, 5'd3};
    assign wire3132 = {5'd5, 5'd3};
    assign wire3133 = {5'd5, 5'd3};
    assign wire3134 = {5'd5, 5'd3};
    assign wire3135 = {5'd5, 5'd3};
    assign wire3136 = {5'd7, 5'd3};
    assign wire3137 = {5'd7, 5'd3};
    assign wire3138 = {5'd7, 5'd3};
    assign wire3139 = {5'd7, 5'd3};
    assign wire3140 = {5'd7, 5'd3};
    assign wire3141 = {5'd7, 5'd3};
    assign wire3142 = {5'd7, 5'd3};
    assign wire3143 = {5'd7, 5'd3};
    assign wire3144 = {5'd7, 5'd3};
    assign wire3145 = {5'd7, 5'd3};
    assign wire3146 = {5'd7, 5'd3};
    assign wire3147 = {5'd7, 5'd3};
    assign wire3148 = {5'd7, 5'd3};
    assign wire3149 = {5'd7, 5'd3};
    assign wire3150 = {5'd7, 5'd3};
    assign wire3151 = {5'd7, 5'd3};
    assign wire3152 = {5'd7, 5'd3};
    assign wire3153 = {5'd7, 5'd3};
    assign wire3154 = {5'd7, 5'd3};
    assign wire3155 = {5'd7, 5'd3};
    assign wire3156 = {5'd7, 5'd3};
    assign wire3157 = {5'd7, 5'd3};
    assign wire3158 = {5'd7, 5'd3};
    assign wire3159 = {5'd7, 5'd3};
    assign wire3160 = {5'd7, 5'd3};
    assign wire3161 = {5'd7, 5'd3};
    assign wire3162 = {5'd7, 5'd3};
    assign wire3163 = {5'd7, 5'd3};
    assign wire3164 = {5'd7, 5'd3};
    assign wire3165 = {5'd7, 5'd3};
    assign wire3166 = {5'd7, 5'd3};
    assign wire3167 = {5'd7, 5'd3};
    assign wire3168 = {5'd9, 5'd3};
    assign wire3169 = {5'd9, 5'd3};
    assign wire3170 = {5'd9, 5'd3};
    assign wire3171 = {5'd9, 5'd3};
    assign wire3172 = {5'd9, 5'd3};
    assign wire3173 = {5'd9, 5'd3};
    assign wire3174 = {5'd9, 5'd3};
    assign wire3175 = {5'd9, 5'd3};
    assign wire3176 = {5'd9, 5'd3};
    assign wire3177 = {5'd9, 5'd3};
    assign wire3178 = {5'd9, 5'd3};
    assign wire3179 = {5'd9, 5'd3};
    assign wire3180 = {5'd9, 5'd3};
    assign wire3181 = {5'd9, 5'd3};
    assign wire3182 = {5'd9, 5'd3};
    assign wire3183 = {5'd9, 5'd3};
    assign wire3184 = {5'd9, 5'd3};
    assign wire3185 = {5'd9, 5'd3};
    assign wire3186 = {5'd9, 5'd3};
    assign wire3187 = {5'd9, 5'd3};
    assign wire3188 = {5'd9, 5'd3};
    assign wire3189 = {5'd9, 5'd3};
    assign wire3190 = {5'd9, 5'd3};
    assign wire3191 = {5'd9, 5'd3};
    assign wire3192 = {5'd9, 5'd3};
    assign wire3193 = {5'd9, 5'd3};
    assign wire3194 = {5'd9, 5'd3};
    assign wire3195 = {5'd9, 5'd3};
    assign wire3196 = {5'd9, 5'd3};
    assign wire3197 = {5'd9, 5'd3};
    assign wire3198 = {5'd9, 5'd3};
    assign wire3199 = {5'd9, 5'd3};
    assign wire3200 = {5'd5, 5'd4};
    assign wire3201 = {5'd5, 5'd4};
    assign wire3202 = {5'd5, 5'd4};
    assign wire3203 = {5'd5, 5'd4};
    assign wire3204 = {5'd6, 5'd5};
    assign wire3205 = {5'd9, 5'd8};
    assign wire3206 = {5'd5, 5'd4};
    assign wire3207 = {5'd5, 5'd4};
    assign wire3208 = {5'd6, 5'd5};
    assign wire3209 = {5'd6, 5'd5};
    assign wire3210 = {5'd6, 5'd5};
    assign wire3211 = {5'd6, 5'd5};
    assign wire3212 = {5'd7, 5'd6};
    assign wire3213 = {5'd6, 5'd5};
    assign wire3214 = {5'd6, 5'd5};
    assign wire3215 = {5'd6, 5'd5};
    assign wire3216 = {5'd9, 5'd8};
    assign wire3217 = {5'd9, 5'd8};
    assign wire3218 = {5'd9, 5'd8};
    assign wire3219 = {5'd9, 5'd8};
    assign wire3220 = {5'd10, 5'd9};
    assign wire3221 = {5'd9, 5'd8};
    assign wire3222 = {5'd9, 5'd8};
    assign wire3223 = {5'd9, 5'd8};
    assign wire3224 = {5'd5, 5'd4};
    assign wire3225 = {5'd5, 5'd4};
    assign wire3226 = {5'd5, 5'd4};
    assign wire3227 = {5'd5, 5'd4};
    assign wire3228 = {5'd5, 5'd4};
    assign wire3229 = {5'd5, 5'd4};
    assign wire3230 = {5'd5, 5'd4};
    assign wire3231 = {5'd5, 5'd4};
    assign wire3232 = {5'd6, 5'd4};
    assign wire3233 = {5'd6, 5'd4};
    assign wire3234 = {5'd6, 5'd4};
    assign wire3235 = {5'd6, 5'd4};
    assign wire3236 = {5'd7, 5'd5};
    assign wire3237 = {5'd10, 5'd8};
    assign wire3238 = {5'd6, 5'd4};
    assign wire3239 = {5'd6, 5'd4};
    assign wire3240 = {5'd7, 5'd5};
    assign wire3241 = {5'd7, 5'd5};
    assign wire3242 = {5'd7, 5'd5};
    assign wire3243 = {5'd7, 5'd5};
    assign wire3244 = {5'd8, 5'd6};
    assign wire3245 = {5'd7, 5'd5};
    assign wire3246 = {5'd7, 5'd5};
    assign wire3247 = {5'd7, 5'd5};
    assign wire3248 = {5'd10, 5'd8};
    assign wire3249 = {5'd10, 5'd8};
    assign wire3250 = {5'd10, 5'd8};
    assign wire3251 = {5'd10, 5'd8};
    assign wire3252 = {5'd11, 5'd9};
    assign wire3253 = {5'd10, 5'd8};
    assign wire3254 = {5'd10, 5'd8};
    assign wire3255 = {5'd10, 5'd8};
    assign wire3256 = {5'd6, 5'd4};
    assign wire3257 = {5'd6, 5'd4};
    assign wire3258 = {5'd6, 5'd4};
    assign wire3259 = {5'd6, 5'd4};
    assign wire3260 = {5'd6, 5'd4};
    assign wire3261 = {5'd6, 5'd4};
    assign wire3262 = {5'd6, 5'd4};
    assign wire3263 = {5'd6, 5'd4};
    assign wire3264 = {5'd8, 5'd4};
    assign wire3265 = {5'd8, 5'd4};
    assign wire3266 = {5'd8, 5'd4};
    assign wire3267 = {5'd8, 5'd4};
    assign wire3268 = {5'd9, 5'd5};
    assign wire3269 = {5'd12, 5'd8};
    assign wire3270 = {5'd8, 5'd4};
    assign wire3271 = {5'd8, 5'd4};
    assign wire3272 = {5'd9, 5'd5};
    assign wire3273 = {5'd9, 5'd5};
    assign wire3274 = {5'd9, 5'd5};
    assign wire3275 = {5'd9, 5'd5};
    assign wire3276 = {5'd10, 5'd6};
    assign wire3277 = {5'd9, 5'd5};
    assign wire3278 = {5'd9, 5'd5};
    assign wire3279 = {5'd9, 5'd5};
    assign wire3280 = {5'd12, 5'd8};
    assign wire3281 = {5'd12, 5'd8};
    assign wire3282 = {5'd12, 5'd8};
    assign wire3283 = {5'd12, 5'd8};
    assign wire3284 = {5'd13, 5'd9};
    assign wire3285 = {5'd12, 5'd8};
    assign wire3286 = {5'd12, 5'd8};
    assign wire3287 = {5'd12, 5'd8};
    assign wire3288 = {5'd8, 5'd4};
    assign wire3289 = {5'd8, 5'd4};
    assign wire3290 = {5'd8, 5'd4};
    assign wire3291 = {5'd8, 5'd4};
    assign wire3292 = {5'd8, 5'd4};
    assign wire3293 = {5'd8, 5'd4};
    assign wire3294 = {5'd8, 5'd4};
    assign wire3295 = {5'd8, 5'd4};
    assign wire3296 = {5'd10, 5'd4};
    assign wire3297 = {5'd10, 5'd4};
    assign wire3298 = {5'd10, 5'd4};
    assign wire3299 = {5'd10, 5'd4};
    assign wire3300 = {5'd11, 5'd5};
    assign wire3301 = {5'd14, 5'd8};
    assign wire3302 = {5'd10, 5'd4};
    assign wire3303 = {5'd10, 5'd4};
    assign wire3304 = {5'd11, 5'd5};
    assign wire3305 = {5'd11, 5'd5};
    assign wire3306 = {5'd11, 5'd5};
    assign wire3307 = {5'd11, 5'd5};
    assign wire3308 = {5'd12, 5'd6};
    assign wire3309 = {5'd11, 5'd5};
    assign wire3310 = {5'd11, 5'd5};
    assign wire3311 = {5'd11, 5'd5};
    assign wire3312 = {5'd14, 5'd8};
    assign wire3313 = {5'd14, 5'd8};
    assign wire3314 = {5'd14, 5'd8};
    assign wire3315 = {5'd14, 5'd8};
    assign wire3316 = {5'd15, 5'd9};
    assign wire3317 = {5'd14, 5'd8};
    assign wire3318 = {5'd14, 5'd8};
    assign wire3319 = {5'd14, 5'd8};
    assign wire3320 = {5'd10, 5'd4};
    assign wire3321 = {5'd10, 5'd4};
    assign wire3322 = {5'd10, 5'd4};
    assign wire3323 = {5'd10, 5'd4};
    assign wire3324 = {5'd10, 5'd4};
    assign wire3325 = {5'd10, 5'd4};
    assign wire3326 = {5'd10, 5'd4};
    assign wire3327 = {5'd10, 5'd4};
    assign wire3328 = {5'd5, 5'd4};
    assign wire3329 = {5'd5, 5'd4};
    assign wire3330 = {5'd5, 5'd4};
    assign wire3331 = {5'd5, 5'd4};
    assign wire3332 = {5'd5, 5'd4};
    assign wire3333 = {5'd5, 5'd4};
    assign wire3334 = {5'd5, 5'd4};
    assign wire3335 = {5'd5, 5'd4};
    assign wire3336 = {5'd5, 5'd4};
    assign wire3337 = {5'd5, 5'd4};
    assign wire3338 = {5'd5, 5'd4};
    assign wire3339 = {5'd5, 5'd4};
    assign wire3340 = {5'd5, 5'd4};
    assign wire3341 = {5'd5, 5'd4};
    assign wire3342 = {5'd5, 5'd4};
    assign wire3343 = {5'd5, 5'd4};
    assign wire3344 = {5'd5, 5'd4};
    assign wire3345 = {5'd5, 5'd4};
    assign wire3346 = {5'd5, 5'd4};
    assign wire3347 = {5'd5, 5'd4};
    assign wire3348 = {5'd5, 5'd4};
    assign wire3349 = {5'd5, 5'd4};
    assign wire3350 = {5'd5, 5'd4};
    assign wire3351 = {5'd5, 5'd4};
    assign wire3352 = {5'd5, 5'd4};
    assign wire3353 = {5'd5, 5'd4};
    assign wire3354 = {5'd5, 5'd4};
    assign wire3355 = {5'd5, 5'd4};
    assign wire3356 = {5'd5, 5'd4};
    assign wire3357 = {5'd5, 5'd4};
    assign wire3358 = {5'd5, 5'd4};
    assign wire3359 = {5'd5, 5'd4};
    assign wire3360 = {5'd6, 5'd4};
    assign wire3361 = {5'd6, 5'd4};
    assign wire3362 = {5'd6, 5'd4};
    assign wire3363 = {5'd6, 5'd4};
    assign wire3364 = {5'd6, 5'd4};
    assign wire3365 = {5'd6, 5'd4};
    assign wire3366 = {5'd6, 5'd4};
    assign wire3367 = {5'd6, 5'd4};
    assign wire3368 = {5'd6, 5'd4};
    assign wire3369 = {5'd6, 5'd4};
    assign wire3370 = {5'd6, 5'd4};
    assign wire3371 = {5'd6, 5'd4};
    assign wire3372 = {5'd6, 5'd4};
    assign wire3373 = {5'd6, 5'd4};
    assign wire3374 = {5'd6, 5'd4};
    assign wire3375 = {5'd6, 5'd4};
    assign wire3376 = {5'd6, 5'd4};
    assign wire3377 = {5'd6, 5'd4};
    assign wire3378 = {5'd6, 5'd4};
    assign wire3379 = {5'd6, 5'd4};
    assign wire3380 = {5'd6, 5'd4};
    assign wire3381 = {5'd6, 5'd4};
    assign wire3382 = {5'd6, 5'd4};
    assign wire3383 = {5'd6, 5'd4};
    assign wire3384 = {5'd6, 5'd4};
    assign wire3385 = {5'd6, 5'd4};
    assign wire3386 = {5'd6, 5'd4};
    assign wire3387 = {5'd6, 5'd4};
    assign wire3388 = {5'd6, 5'd4};
    assign wire3389 = {5'd6, 5'd4};
    assign wire3390 = {5'd6, 5'd4};
    assign wire3391 = {5'd6, 5'd4};
    assign wire3392 = {5'd8, 5'd4};
    assign wire3393 = {5'd8, 5'd4};
    assign wire3394 = {5'd8, 5'd4};
    assign wire3395 = {5'd8, 5'd4};
    assign wire3396 = {5'd8, 5'd4};
    assign wire3397 = {5'd8, 5'd4};
    assign wire3398 = {5'd8, 5'd4};
    assign wire3399 = {5'd8, 5'd4};
    assign wire3400 = {5'd8, 5'd4};
    assign wire3401 = {5'd8, 5'd4};
    assign wire3402 = {5'd8, 5'd4};
    assign wire3403 = {5'd8, 5'd4};
    assign wire3404 = {5'd8, 5'd4};
    assign wire3405 = {5'd8, 5'd4};
    assign wire3406 = {5'd8, 5'd4};
    assign wire3407 = {5'd8, 5'd4};
    assign wire3408 = {5'd8, 5'd4};
    assign wire3409 = {5'd8, 5'd4};
    assign wire3410 = {5'd8, 5'd4};
    assign wire3411 = {5'd8, 5'd4};
    assign wire3412 = {5'd8, 5'd4};
    assign wire3413 = {5'd8, 5'd4};
    assign wire3414 = {5'd8, 5'd4};
    assign wire3415 = {5'd8, 5'd4};
    assign wire3416 = {5'd8, 5'd4};
    assign wire3417 = {5'd8, 5'd4};
    assign wire3418 = {5'd8, 5'd4};
    assign wire3419 = {5'd8, 5'd4};
    assign wire3420 = {5'd8, 5'd4};
    assign wire3421 = {5'd8, 5'd4};
    assign wire3422 = {5'd8, 5'd4};
    assign wire3423 = {5'd8, 5'd4};
    assign wire3424 = {5'd10, 5'd4};
    assign wire3425 = {5'd10, 5'd4};
    assign wire3426 = {5'd10, 5'd4};
    assign wire3427 = {5'd10, 5'd4};
    assign wire3428 = {5'd10, 5'd4};
    assign wire3429 = {5'd10, 5'd4};
    assign wire3430 = {5'd10, 5'd4};
    assign wire3431 = {5'd10, 5'd4};
    assign wire3432 = {5'd10, 5'd4};
    assign wire3433 = {5'd10, 5'd4};
    assign wire3434 = {5'd10, 5'd4};
    assign wire3435 = {5'd10, 5'd4};
    assign wire3436 = {5'd10, 5'd4};
    assign wire3437 = {5'd10, 5'd4};
    assign wire3438 = {5'd10, 5'd4};
    assign wire3439 = {5'd10, 5'd4};
    assign wire3440 = {5'd10, 5'd4};
    assign wire3441 = {5'd10, 5'd4};
    assign wire3442 = {5'd10, 5'd4};
    assign wire3443 = {5'd10, 5'd4};
    assign wire3444 = {5'd10, 5'd4};
    assign wire3445 = {5'd10, 5'd4};
    assign wire3446 = {5'd10, 5'd4};
    assign wire3447 = {5'd10, 5'd4};
    assign wire3448 = {5'd10, 5'd4};
    assign wire3449 = {5'd10, 5'd4};
    assign wire3450 = {5'd10, 5'd4};
    assign wire3451 = {5'd10, 5'd4};
    assign wire3452 = {5'd10, 5'd4};
    assign wire3453 = {5'd10, 5'd4};
    assign wire3454 = {5'd10, 5'd4};
    assign wire3455 = {5'd10, 5'd4};
    assign wire3456 = {5'd6, 5'd5};
    assign wire3457 = {5'd6, 5'd5};
    assign wire3458 = {5'd6, 5'd5};
    assign wire3459 = {5'd6, 5'd5};
    assign wire3460 = {5'd7, 5'd6};
    assign wire3461 = {5'd10, 5'd9};
    assign wire3462 = {5'd6, 5'd5};
    assign wire3463 = {5'd6, 5'd5};
    assign wire3464 = {5'd7, 5'd6};
    assign wire3465 = {5'd7, 5'd6};
    assign wire3466 = {5'd7, 5'd6};
    assign wire3467 = {5'd7, 5'd6};
    assign wire3468 = {5'd8, 5'd7};
    assign wire3469 = {5'd7, 5'd6};
    assign wire3470 = {5'd7, 5'd6};
    assign wire3471 = {5'd7, 5'd6};
    assign wire3472 = {5'd10, 5'd9};
    assign wire3473 = {5'd10, 5'd9};
    assign wire3474 = {5'd10, 5'd9};
    assign wire3475 = {5'd10, 5'd9};
    assign wire3476 = {5'd11, 5'd10};
    assign wire3477 = {5'd10, 5'd9};
    assign wire3478 = {5'd10, 5'd9};
    assign wire3479 = {5'd10, 5'd9};
    assign wire3480 = {5'd6, 5'd5};
    assign wire3481 = {5'd6, 5'd5};
    assign wire3482 = {5'd6, 5'd5};
    assign wire3483 = {5'd6, 5'd5};
    assign wire3484 = {5'd6, 5'd5};
    assign wire3485 = {5'd6, 5'd5};
    assign wire3486 = {5'd6, 5'd5};
    assign wire3487 = {5'd6, 5'd5};
    assign wire3488 = {5'd7, 5'd5};
    assign wire3489 = {5'd7, 5'd5};
    assign wire3490 = {5'd7, 5'd5};
    assign wire3491 = {5'd7, 5'd5};
    assign wire3492 = {5'd8, 5'd6};
    assign wire3493 = {5'd11, 5'd9};
    assign wire3494 = {5'd7, 5'd5};
    assign wire3495 = {5'd7, 5'd5};
    assign wire3496 = {5'd8, 5'd6};
    assign wire3497 = {5'd8, 5'd6};
    assign wire3498 = {5'd8, 5'd6};
    assign wire3499 = {5'd8, 5'd6};
    assign wire3500 = {5'd9, 5'd7};
    assign wire3501 = {5'd8, 5'd6};
    assign wire3502 = {5'd8, 5'd6};
    assign wire3503 = {5'd8, 5'd6};
    assign wire3504 = {5'd11, 5'd9};
    assign wire3505 = {5'd11, 5'd9};
    assign wire3506 = {5'd11, 5'd9};
    assign wire3507 = {5'd11, 5'd9};
    assign wire3508 = {5'd12, 5'd10};
    assign wire3509 = {5'd11, 5'd9};
    assign wire3510 = {5'd11, 5'd9};
    assign wire3511 = {5'd11, 5'd9};
    assign wire3512 = {5'd7, 5'd5};
    assign wire3513 = {5'd7, 5'd5};
    assign wire3514 = {5'd7, 5'd5};
    assign wire3515 = {5'd7, 5'd5};
    assign wire3516 = {5'd7, 5'd5};
    assign wire3517 = {5'd7, 5'd5};
    assign wire3518 = {5'd7, 5'd5};
    assign wire3519 = {5'd7, 5'd5};
    assign wire3520 = {5'd9, 5'd5};
    assign wire3521 = {5'd9, 5'd5};
    assign wire3522 = {5'd9, 5'd5};
    assign wire3523 = {5'd9, 5'd5};
    assign wire3524 = {5'd10, 5'd6};
    assign wire3525 = {5'd13, 5'd9};
    assign wire3526 = {5'd9, 5'd5};
    assign wire3527 = {5'd9, 5'd5};
    assign wire3528 = {5'd10, 5'd6};
    assign wire3529 = {5'd10, 5'd6};
    assign wire3530 = {5'd10, 5'd6};
    assign wire3531 = {5'd10, 5'd6};
    assign wire3532 = {5'd11, 5'd7};
    assign wire3533 = {5'd10, 5'd6};
    assign wire3534 = {5'd10, 5'd6};
    assign wire3535 = {5'd10, 5'd6};
    assign wire3536 = {5'd13, 5'd9};
    assign wire3537 = {5'd13, 5'd9};
    assign wire3538 = {5'd13, 5'd9};
    assign wire3539 = {5'd13, 5'd9};
    assign wire3540 = {5'd14, 5'd10};
    assign wire3541 = {5'd13, 5'd9};
    assign wire3542 = {5'd13, 5'd9};
    assign wire3543 = {5'd13, 5'd9};
    assign wire3544 = {5'd9, 5'd5};
    assign wire3545 = {5'd9, 5'd5};
    assign wire3546 = {5'd9, 5'd5};
    assign wire3547 = {5'd9, 5'd5};
    assign wire3548 = {5'd9, 5'd5};
    assign wire3549 = {5'd9, 5'd5};
    assign wire3550 = {5'd9, 5'd5};
    assign wire3551 = {5'd9, 5'd5};
    assign wire3552 = {5'd11, 5'd5};
    assign wire3553 = {5'd11, 5'd5};
    assign wire3554 = {5'd11, 5'd5};
    assign wire3555 = {5'd11, 5'd5};
    assign wire3556 = {5'd12, 5'd6};
    assign wire3557 = {5'd15, 5'd9};
    assign wire3558 = {5'd11, 5'd5};
    assign wire3559 = {5'd11, 5'd5};
    assign wire3560 = {5'd12, 5'd6};
    assign wire3561 = {5'd12, 5'd6};
    assign wire3562 = {5'd12, 5'd6};
    assign wire3563 = {5'd12, 5'd6};
    assign wire3564 = {5'd13, 5'd7};
    assign wire3565 = {5'd12, 5'd6};
    assign wire3566 = {5'd12, 5'd6};
    assign wire3567 = {5'd12, 5'd6};
    assign wire3568 = {5'd15, 5'd9};
    assign wire3569 = {5'd15, 5'd9};
    assign wire3570 = {5'd15, 5'd9};
    assign wire3571 = {5'd15, 5'd9};
    assign wire3572 = {5'd16, 5'd10};
    assign wire3573 = {5'd15, 5'd9};
    assign wire3574 = {5'd15, 5'd9};
    assign wire3575 = {5'd15, 5'd9};
    assign wire3576 = {5'd11, 5'd5};
    assign wire3577 = {5'd11, 5'd5};
    assign wire3578 = {5'd11, 5'd5};
    assign wire3579 = {5'd11, 5'd5};
    assign wire3580 = {5'd11, 5'd5};
    assign wire3581 = {5'd11, 5'd5};
    assign wire3582 = {5'd11, 5'd5};
    assign wire3583 = {5'd11, 5'd5};
    assign wire3584 = {5'd5, 5'd4};
    assign wire3585 = {5'd5, 5'd4};
    assign wire3586 = {5'd5, 5'd4};
    assign wire3587 = {5'd5, 5'd4};
    assign wire3588 = {5'd5, 5'd4};
    assign wire3589 = {5'd5, 5'd4};
    assign wire3590 = {5'd5, 5'd4};
    assign wire3591 = {5'd5, 5'd4};
    assign wire3592 = {5'd5, 5'd4};
    assign wire3593 = {5'd5, 5'd4};
    assign wire3594 = {5'd5, 5'd4};
    assign wire3595 = {5'd5, 5'd4};
    assign wire3596 = {5'd5, 5'd4};
    assign wire3597 = {5'd5, 5'd4};
    assign wire3598 = {5'd5, 5'd4};
    assign wire3599 = {5'd5, 5'd4};
    assign wire3600 = {5'd5, 5'd4};
    assign wire3601 = {5'd5, 5'd4};
    assign wire3602 = {5'd5, 5'd4};
    assign wire3603 = {5'd5, 5'd4};
    assign wire3604 = {5'd5, 5'd4};
    assign wire3605 = {5'd5, 5'd4};
    assign wire3606 = {5'd5, 5'd4};
    assign wire3607 = {5'd5, 5'd4};
    assign wire3608 = {5'd5, 5'd4};
    assign wire3609 = {5'd5, 5'd4};
    assign wire3610 = {5'd5, 5'd4};
    assign wire3611 = {5'd5, 5'd4};
    assign wire3612 = {5'd5, 5'd4};
    assign wire3613 = {5'd5, 5'd4};
    assign wire3614 = {5'd5, 5'd4};
    assign wire3615 = {5'd5, 5'd4};
    assign wire3616 = {5'd6, 5'd4};
    assign wire3617 = {5'd6, 5'd4};
    assign wire3618 = {5'd6, 5'd4};
    assign wire3619 = {5'd6, 5'd4};
    assign wire3620 = {5'd6, 5'd4};
    assign wire3621 = {5'd6, 5'd4};
    assign wire3622 = {5'd6, 5'd4};
    assign wire3623 = {5'd6, 5'd4};
    assign wire3624 = {5'd6, 5'd4};
    assign wire3625 = {5'd6, 5'd4};
    assign wire3626 = {5'd6, 5'd4};
    assign wire3627 = {5'd6, 5'd4};
    assign wire3628 = {5'd6, 5'd4};
    assign wire3629 = {5'd6, 5'd4};
    assign wire3630 = {5'd6, 5'd4};
    assign wire3631 = {5'd6, 5'd4};
    assign wire3632 = {5'd6, 5'd4};
    assign wire3633 = {5'd6, 5'd4};
    assign wire3634 = {5'd6, 5'd4};
    assign wire3635 = {5'd6, 5'd4};
    assign wire3636 = {5'd6, 5'd4};
    assign wire3637 = {5'd6, 5'd4};
    assign wire3638 = {5'd6, 5'd4};
    assign wire3639 = {5'd6, 5'd4};
    assign wire3640 = {5'd6, 5'd4};
    assign wire3641 = {5'd6, 5'd4};
    assign wire3642 = {5'd6, 5'd4};
    assign wire3643 = {5'd6, 5'd4};
    assign wire3644 = {5'd6, 5'd4};
    assign wire3645 = {5'd6, 5'd4};
    assign wire3646 = {5'd6, 5'd4};
    assign wire3647 = {5'd6, 5'd4};
    assign wire3648 = {5'd8, 5'd4};
    assign wire3649 = {5'd8, 5'd4};
    assign wire3650 = {5'd8, 5'd4};
    assign wire3651 = {5'd8, 5'd4};
    assign wire3652 = {5'd8, 5'd4};
    assign wire3653 = {5'd8, 5'd4};
    assign wire3654 = {5'd8, 5'd4};
    assign wire3655 = {5'd8, 5'd4};
    assign wire3656 = {5'd8, 5'd4};
    assign wire3657 = {5'd8, 5'd4};
    assign wire3658 = {5'd8, 5'd4};
    assign wire3659 = {5'd8, 5'd4};
    assign wire3660 = {5'd8, 5'd4};
    assign wire3661 = {5'd8, 5'd4};
    assign wire3662 = {5'd8, 5'd4};
    assign wire3663 = {5'd8, 5'd4};
    assign wire3664 = {5'd8, 5'd4};
    assign wire3665 = {5'd8, 5'd4};
    assign wire3666 = {5'd8, 5'd4};
    assign wire3667 = {5'd8, 5'd4};
    assign wire3668 = {5'd8, 5'd4};
    assign wire3669 = {5'd8, 5'd4};
    assign wire3670 = {5'd8, 5'd4};
    assign wire3671 = {5'd8, 5'd4};
    assign wire3672 = {5'd8, 5'd4};
    assign wire3673 = {5'd8, 5'd4};
    assign wire3674 = {5'd8, 5'd4};
    assign wire3675 = {5'd8, 5'd4};
    assign wire3676 = {5'd8, 5'd4};
    assign wire3677 = {5'd8, 5'd4};
    assign wire3678 = {5'd8, 5'd4};
    assign wire3679 = {5'd8, 5'd4};
    assign wire3680 = {5'd10, 5'd4};
    assign wire3681 = {5'd10, 5'd4};
    assign wire3682 = {5'd10, 5'd4};
    assign wire3683 = {5'd10, 5'd4};
    assign wire3684 = {5'd10, 5'd4};
    assign wire3685 = {5'd10, 5'd4};
    assign wire3686 = {5'd10, 5'd4};
    assign wire3687 = {5'd10, 5'd4};
    assign wire3688 = {5'd10, 5'd4};
    assign wire3689 = {5'd10, 5'd4};
    assign wire3690 = {5'd10, 5'd4};
    assign wire3691 = {5'd10, 5'd4};
    assign wire3692 = {5'd10, 5'd4};
    assign wire3693 = {5'd10, 5'd4};
    assign wire3694 = {5'd10, 5'd4};
    assign wire3695 = {5'd10, 5'd4};
    assign wire3696 = {5'd10, 5'd4};
    assign wire3697 = {5'd10, 5'd4};
    assign wire3698 = {5'd10, 5'd4};
    assign wire3699 = {5'd10, 5'd4};
    assign wire3700 = {5'd10, 5'd4};
    assign wire3701 = {5'd10, 5'd4};
    assign wire3702 = {5'd10, 5'd4};
    assign wire3703 = {5'd10, 5'd4};
    assign wire3704 = {5'd10, 5'd4};
    assign wire3705 = {5'd10, 5'd4};
    assign wire3706 = {5'd10, 5'd4};
    assign wire3707 = {5'd10, 5'd4};
    assign wire3708 = {5'd10, 5'd4};
    assign wire3709 = {5'd10, 5'd4};
    assign wire3710 = {5'd10, 5'd4};
    assign wire3711 = {5'd10, 5'd4};
    assign wire3712 = {5'd6, 5'd5};
    assign wire3713 = {5'd6, 5'd5};
    assign wire3714 = {5'd6, 5'd5};
    assign wire3715 = {5'd6, 5'd5};
    assign wire3716 = {5'd6, 5'd5};
    assign wire3717 = {5'd8, 5'd7};
    assign wire3718 = {5'd6, 5'd5};
    assign wire3719 = {5'd6, 5'd5};
    assign wire3720 = {5'd7, 5'd6};
    assign wire3721 = {5'd7, 5'd6};
    assign wire3722 = {5'd7, 5'd6};
    assign wire3723 = {5'd7, 5'd6};
    assign wire3724 = {5'd7, 5'd6};
    assign wire3725 = {5'd7, 5'd6};
    assign wire3726 = {5'd7, 5'd6};
    assign wire3727 = {5'd7, 5'd6};
    assign wire3728 = {5'd8, 5'd7};
    assign wire3729 = {5'd8, 5'd7};
    assign wire3730 = {5'd8, 5'd7};
    assign wire3731 = {5'd8, 5'd7};
    assign wire3732 = {5'd8, 5'd7};
    assign wire3733 = {5'd8, 5'd7};
    assign wire3734 = {5'd8, 5'd7};
    assign wire3735 = {5'd8, 5'd7};
    assign wire3736 = {5'd6, 5'd5};
    assign wire3737 = {5'd6, 5'd5};
    assign wire3738 = {5'd6, 5'd5};
    assign wire3739 = {5'd6, 5'd5};
    assign wire3740 = {5'd6, 5'd5};
    assign wire3741 = {5'd6, 5'd5};
    assign wire3742 = {5'd6, 5'd5};
    assign wire3743 = {5'd6, 5'd5};
    assign wire3744 = {5'd7, 5'd5};
    assign wire3745 = {5'd7, 5'd5};
    assign wire3746 = {5'd7, 5'd5};
    assign wire3747 = {5'd7, 5'd5};
    assign wire3748 = {5'd7, 5'd5};
    assign wire3749 = {5'd9, 5'd7};
    assign wire3750 = {5'd7, 5'd5};
    assign wire3751 = {5'd7, 5'd5};
    assign wire3752 = {5'd8, 5'd6};
    assign wire3753 = {5'd8, 5'd6};
    assign wire3754 = {5'd8, 5'd6};
    assign wire3755 = {5'd8, 5'd6};
    assign wire3756 = {5'd8, 5'd6};
    assign wire3757 = {5'd8, 5'd6};
    assign wire3758 = {5'd8, 5'd6};
    assign wire3759 = {5'd8, 5'd6};
    assign wire3760 = {5'd9, 5'd7};
    assign wire3761 = {5'd9, 5'd7};
    assign wire3762 = {5'd9, 5'd7};
    assign wire3763 = {5'd9, 5'd7};
    assign wire3764 = {5'd9, 5'd7};
    assign wire3765 = {5'd9, 5'd7};
    assign wire3766 = {5'd9, 5'd7};
    assign wire3767 = {5'd9, 5'd7};
    assign wire3768 = {5'd7, 5'd5};
    assign wire3769 = {5'd7, 5'd5};
    assign wire3770 = {5'd7, 5'd5};
    assign wire3771 = {5'd7, 5'd5};
    assign wire3772 = {5'd7, 5'd5};
    assign wire3773 = {5'd7, 5'd5};
    assign wire3774 = {5'd7, 5'd5};
    assign wire3775 = {5'd7, 5'd5};
    assign wire3776 = {5'd9, 5'd5};
    assign wire3777 = {5'd9, 5'd5};
    assign wire3778 = {5'd9, 5'd5};
    assign wire3779 = {5'd9, 5'd5};
    assign wire3780 = {5'd9, 5'd5};
    assign wire3781 = {5'd11, 5'd7};
    assign wire3782 = {5'd9, 5'd5};
    assign wire3783 = {5'd9, 5'd5};
    assign wire3784 = {5'd10, 5'd6};
    assign wire3785 = {5'd10, 5'd6};
    assign wire3786 = {5'd10, 5'd6};
    assign wire3787 = {5'd10, 5'd6};
    assign wire3788 = {5'd10, 5'd6};
    assign wire3789 = {5'd10, 5'd6};
    assign wire3790 = {5'd10, 5'd6};
    assign wire3791 = {5'd10, 5'd6};
    assign wire3792 = {5'd11, 5'd7};
    assign wire3793 = {5'd11, 5'd7};
    assign wire3794 = {5'd11, 5'd7};
    assign wire3795 = {5'd11, 5'd7};
    assign wire3796 = {5'd11, 5'd7};
    assign wire3797 = {5'd11, 5'd7};
    assign wire3798 = {5'd11, 5'd7};
    assign wire3799 = {5'd11, 5'd7};
    assign wire3800 = {5'd9, 5'd5};
    assign wire3801 = {5'd9, 5'd5};
    assign wire3802 = {5'd9, 5'd5};
    assign wire3803 = {5'd9, 5'd5};
    assign wire3804 = {5'd9, 5'd5};
    assign wire3805 = {5'd9, 5'd5};
    assign wire3806 = {5'd9, 5'd5};
    assign wire3807 = {5'd9, 5'd5};
    assign wire3808 = {5'd11, 5'd5};
    assign wire3809 = {5'd11, 5'd5};
    assign wire3810 = {5'd11, 5'd5};
    assign wire3811 = {5'd11, 5'd5};
    assign wire3812 = {5'd11, 5'd5};
    assign wire3813 = {5'd13, 5'd7};
    assign wire3814 = {5'd11, 5'd5};
    assign wire3815 = {5'd11, 5'd5};
    assign wire3816 = {5'd12, 5'd6};
    assign wire3817 = {5'd12, 5'd6};
    assign wire3818 = {5'd12, 5'd6};
    assign wire3819 = {5'd12, 5'd6};
    assign wire3820 = {5'd12, 5'd6};
    assign wire3821 = {5'd12, 5'd6};
    assign wire3822 = {5'd12, 5'd6};
    assign wire3823 = {5'd12, 5'd6};
    assign wire3824 = {5'd13, 5'd7};
    assign wire3825 = {5'd13, 5'd7};
    assign wire3826 = {5'd13, 5'd7};
    assign wire3827 = {5'd13, 5'd7};
    assign wire3828 = {5'd13, 5'd7};
    assign wire3829 = {5'd13, 5'd7};
    assign wire3830 = {5'd13, 5'd7};
    assign wire3831 = {5'd13, 5'd7};
    assign wire3832 = {5'd11, 5'd5};
    assign wire3833 = {5'd11, 5'd5};
    assign wire3834 = {5'd11, 5'd5};
    assign wire3835 = {5'd11, 5'd5};
    assign wire3836 = {5'd11, 5'd5};
    assign wire3837 = {5'd11, 5'd5};
    assign wire3838 = {5'd11, 5'd5};
    assign wire3839 = {5'd11, 5'd5};
    assign wire3840 = {5'd6, 5'd5};
    assign wire3841 = {5'd6, 5'd5};
    assign wire3842 = {5'd6, 5'd5};
    assign wire3843 = {5'd6, 5'd5};
    assign wire3844 = {5'd6, 5'd5};
    assign wire3845 = {5'd6, 5'd5};
    assign wire3846 = {5'd6, 5'd5};
    assign wire3847 = {5'd6, 5'd5};
    assign wire3848 = {5'd6, 5'd5};
    assign wire3849 = {5'd6, 5'd5};
    assign wire3850 = {5'd6, 5'd5};
    assign wire3851 = {5'd6, 5'd5};
    assign wire3852 = {5'd6, 5'd5};
    assign wire3853 = {5'd6, 5'd5};
    assign wire3854 = {5'd6, 5'd5};
    assign wire3855 = {5'd6, 5'd5};
    assign wire3856 = {5'd6, 5'd5};
    assign wire3857 = {5'd6, 5'd5};
    assign wire3858 = {5'd6, 5'd5};
    assign wire3859 = {5'd6, 5'd5};
    assign wire3860 = {5'd6, 5'd5};
    assign wire3861 = {5'd6, 5'd5};
    assign wire3862 = {5'd6, 5'd5};
    assign wire3863 = {5'd6, 5'd5};
    assign wire3864 = {5'd6, 5'd5};
    assign wire3865 = {5'd6, 5'd5};
    assign wire3866 = {5'd6, 5'd5};
    assign wire3867 = {5'd6, 5'd5};
    assign wire3868 = {5'd6, 5'd5};
    assign wire3869 = {5'd6, 5'd5};
    assign wire3870 = {5'd6, 5'd5};
    assign wire3871 = {5'd6, 5'd5};
    assign wire3872 = {5'd7, 5'd5};
    assign wire3873 = {5'd7, 5'd5};
    assign wire3874 = {5'd7, 5'd5};
    assign wire3875 = {5'd7, 5'd5};
    assign wire3876 = {5'd7, 5'd5};
    assign wire3877 = {5'd7, 5'd5};
    assign wire3878 = {5'd7, 5'd5};
    assign wire3879 = {5'd7, 5'd5};
    assign wire3880 = {5'd7, 5'd5};
    assign wire3881 = {5'd7, 5'd5};
    assign wire3882 = {5'd7, 5'd5};
    assign wire3883 = {5'd7, 5'd5};
    assign wire3884 = {5'd7, 5'd5};
    assign wire3885 = {5'd7, 5'd5};
    assign wire3886 = {5'd7, 5'd5};
    assign wire3887 = {5'd7, 5'd5};
    assign wire3888 = {5'd7, 5'd5};
    assign wire3889 = {5'd7, 5'd5};
    assign wire3890 = {5'd7, 5'd5};
    assign wire3891 = {5'd7, 5'd5};
    assign wire3892 = {5'd7, 5'd5};
    assign wire3893 = {5'd7, 5'd5};
    assign wire3894 = {5'd7, 5'd5};
    assign wire3895 = {5'd7, 5'd5};
    assign wire3896 = {5'd7, 5'd5};
    assign wire3897 = {5'd7, 5'd5};
    assign wire3898 = {5'd7, 5'd5};
    assign wire3899 = {5'd7, 5'd5};
    assign wire3900 = {5'd7, 5'd5};
    assign wire3901 = {5'd7, 5'd5};
    assign wire3902 = {5'd7, 5'd5};
    assign wire3903 = {5'd7, 5'd5};
    assign wire3904 = {5'd9, 5'd5};
    assign wire3905 = {5'd9, 5'd5};
    assign wire3906 = {5'd9, 5'd5};
    assign wire3907 = {5'd9, 5'd5};
    assign wire3908 = {5'd9, 5'd5};
    assign wire3909 = {5'd9, 5'd5};
    assign wire3910 = {5'd9, 5'd5};
    assign wire3911 = {5'd9, 5'd5};
    assign wire3912 = {5'd9, 5'd5};
    assign wire3913 = {5'd9, 5'd5};
    assign wire3914 = {5'd9, 5'd5};
    assign wire3915 = {5'd9, 5'd5};
    assign wire3916 = {5'd9, 5'd5};
    assign wire3917 = {5'd9, 5'd5};
    assign wire3918 = {5'd9, 5'd5};
    assign wire3919 = {5'd9, 5'd5};
    assign wire3920 = {5'd9, 5'd5};
    assign wire3921 = {5'd9, 5'd5};
    assign wire3922 = {5'd9, 5'd5};
    assign wire3923 = {5'd9, 5'd5};
    assign wire3924 = {5'd9, 5'd5};
    assign wire3925 = {5'd9, 5'd5};
    assign wire3926 = {5'd9, 5'd5};
    assign wire3927 = {5'd9, 5'd5};
    assign wire3928 = {5'd9, 5'd5};
    assign wire3929 = {5'd9, 5'd5};
    assign wire3930 = {5'd9, 5'd5};
    assign wire3931 = {5'd9, 5'd5};
    assign wire3932 = {5'd9, 5'd5};
    assign wire3933 = {5'd9, 5'd5};
    assign wire3934 = {5'd9, 5'd5};
    assign wire3935 = {5'd9, 5'd5};
    assign wire3936 = {5'd11, 5'd5};
    assign wire3937 = {5'd11, 5'd5};
    assign wire3938 = {5'd11, 5'd5};
    assign wire3939 = {5'd11, 5'd5};
    assign wire3940 = {5'd11, 5'd5};
    assign wire3941 = {5'd11, 5'd5};
    assign wire3942 = {5'd11, 5'd5};
    assign wire3943 = {5'd11, 5'd5};
    assign wire3944 = {5'd11, 5'd5};
    assign wire3945 = {5'd11, 5'd5};
    assign wire3946 = {5'd11, 5'd5};
    assign wire3947 = {5'd11, 5'd5};
    assign wire3948 = {5'd11, 5'd5};
    assign wire3949 = {5'd11, 5'd5};
    assign wire3950 = {5'd11, 5'd5};
    assign wire3951 = {5'd11, 5'd5};
    assign wire3952 = {5'd11, 5'd5};
    assign wire3953 = {5'd11, 5'd5};
    assign wire3954 = {5'd11, 5'd5};
    assign wire3955 = {5'd11, 5'd5};
    assign wire3956 = {5'd11, 5'd5};
    assign wire3957 = {5'd11, 5'd5};
    assign wire3958 = {5'd11, 5'd5};
    assign wire3959 = {5'd11, 5'd5};
    assign wire3960 = {5'd11, 5'd5};
    assign wire3961 = {5'd11, 5'd5};
    assign wire3962 = {5'd11, 5'd5};
    assign wire3963 = {5'd11, 5'd5};
    assign wire3964 = {5'd11, 5'd5};
    assign wire3965 = {5'd11, 5'd5};
    assign wire3966 = {5'd11, 5'd5};
    assign wire3967 = {5'd11, 5'd5};
    assign wire3968 = {5'd7, 5'd6};
    assign wire3969 = {5'd7, 5'd6};
    assign wire3970 = {5'd7, 5'd6};
    assign wire3971 = {5'd7, 5'd6};
    assign wire3972 = {5'd7, 5'd6};
    assign wire3973 = {5'd9, 5'd8};
    assign wire3974 = {5'd7, 5'd6};
    assign wire3975 = {5'd7, 5'd6};
    assign wire3976 = {5'd8, 5'd7};
    assign wire3977 = {5'd8, 5'd7};
    assign wire3978 = {5'd8, 5'd7};
    assign wire3979 = {5'd8, 5'd7};
    assign wire3980 = {5'd8, 5'd7};
    assign wire3981 = {5'd8, 5'd7};
    assign wire3982 = {5'd8, 5'd7};
    assign wire3983 = {5'd8, 5'd7};
    assign wire3984 = {5'd9, 5'd8};
    assign wire3985 = {5'd9, 5'd8};
    assign wire3986 = {5'd9, 5'd8};
    assign wire3987 = {5'd9, 5'd8};
    assign wire3988 = {5'd9, 5'd8};
    assign wire3989 = {5'd9, 5'd8};
    assign wire3990 = {5'd9, 5'd8};
    assign wire3991 = {5'd9, 5'd8};
    assign wire3992 = {5'd7, 5'd6};
    assign wire3993 = {5'd7, 5'd6};
    assign wire3994 = {5'd7, 5'd6};
    assign wire3995 = {5'd7, 5'd6};
    assign wire3996 = {5'd7, 5'd6};
    assign wire3997 = {5'd7, 5'd6};
    assign wire3998 = {5'd7, 5'd6};
    assign wire3999 = {5'd7, 5'd6};
    assign wire4000 = {5'd8, 5'd6};
    assign wire4001 = {5'd8, 5'd6};
    assign wire4002 = {5'd8, 5'd6};
    assign wire4003 = {5'd8, 5'd6};
    assign wire4004 = {5'd8, 5'd6};
    assign wire4005 = {5'd10, 5'd8};
    assign wire4006 = {5'd8, 5'd6};
    assign wire4007 = {5'd8, 5'd6};
    assign wire4008 = {5'd9, 5'd7};
    assign wire4009 = {5'd9, 5'd7};
    assign wire4010 = {5'd9, 5'd7};
    assign wire4011 = {5'd9, 5'd7};
    assign wire4012 = {5'd9, 5'd7};
    assign wire4013 = {5'd9, 5'd7};
    assign wire4014 = {5'd9, 5'd7};
    assign wire4015 = {5'd9, 5'd7};
    assign wire4016 = {5'd10, 5'd8};
    assign wire4017 = {5'd10, 5'd8};
    assign wire4018 = {5'd10, 5'd8};
    assign wire4019 = {5'd10, 5'd8};
    assign wire4020 = {5'd10, 5'd8};
    assign wire4021 = {5'd10, 5'd8};
    assign wire4022 = {5'd10, 5'd8};
    assign wire4023 = {5'd10, 5'd8};
    assign wire4024 = {5'd8, 5'd6};
    assign wire4025 = {5'd8, 5'd6};
    assign wire4026 = {5'd8, 5'd6};
    assign wire4027 = {5'd8, 5'd6};
    assign wire4028 = {5'd8, 5'd6};
    assign wire4029 = {5'd8, 5'd6};
    assign wire4030 = {5'd8, 5'd6};
    assign wire4031 = {5'd8, 5'd6};
    assign wire4032 = {5'd10, 5'd6};
    assign wire4033 = {5'd10, 5'd6};
    assign wire4034 = {5'd10, 5'd6};
    assign wire4035 = {5'd10, 5'd6};
    assign wire4036 = {5'd10, 5'd6};
    assign wire4037 = {5'd12, 5'd8};
    assign wire4038 = {5'd10, 5'd6};
    assign wire4039 = {5'd10, 5'd6};
    assign wire4040 = {5'd11, 5'd7};
    assign wire4041 = {5'd11, 5'd7};
    assign wire4042 = {5'd11, 5'd7};
    assign wire4043 = {5'd11, 5'd7};
    assign wire4044 = {5'd11, 5'd7};
    assign wire4045 = {5'd11, 5'd7};
    assign wire4046 = {5'd11, 5'd7};
    assign wire4047 = {5'd11, 5'd7};
    assign wire4048 = {5'd12, 5'd8};
    assign wire4049 = {5'd12, 5'd8};
    assign wire4050 = {5'd12, 5'd8};
    assign wire4051 = {5'd12, 5'd8};
    assign wire4052 = {5'd12, 5'd8};
    assign wire4053 = {5'd12, 5'd8};
    assign wire4054 = {5'd12, 5'd8};
    assign wire4055 = {5'd12, 5'd8};
    assign wire4056 = {5'd10, 5'd6};
    assign wire4057 = {5'd10, 5'd6};
    assign wire4058 = {5'd10, 5'd6};
    assign wire4059 = {5'd10, 5'd6};
    assign wire4060 = {5'd10, 5'd6};
    assign wire4061 = {5'd10, 5'd6};
    assign wire4062 = {5'd10, 5'd6};
    assign wire4063 = {5'd10, 5'd6};
    assign wire4064 = {5'd12, 5'd6};
    assign wire4065 = {5'd12, 5'd6};
    assign wire4066 = {5'd12, 5'd6};
    assign wire4067 = {5'd12, 5'd6};
    assign wire4068 = {5'd12, 5'd6};
    assign wire4069 = {5'd14, 5'd8};
    assign wire4070 = {5'd12, 5'd6};
    assign wire4071 = {5'd12, 5'd6};
    assign wire4072 = {5'd13, 5'd7};
    assign wire4073 = {5'd13, 5'd7};
    assign wire4074 = {5'd13, 5'd7};
    assign wire4075 = {5'd13, 5'd7};
    assign wire4076 = {5'd13, 5'd7};
    assign wire4077 = {5'd13, 5'd7};
    assign wire4078 = {5'd13, 5'd7};
    assign wire4079 = {5'd13, 5'd7};
    assign wire4080 = {5'd14, 5'd8};
    assign wire4081 = {5'd14, 5'd8};
    assign wire4082 = {5'd14, 5'd8};
    assign wire4083 = {5'd14, 5'd8};
    assign wire4084 = {5'd14, 5'd8};
    assign wire4085 = {5'd14, 5'd8};
    assign wire4086 = {5'd14, 5'd8};
    assign wire4087 = {5'd14, 5'd8};
    assign wire4088 = {5'd12, 5'd6};
    assign wire4089 = {5'd12, 5'd6};
    assign wire4090 = {5'd12, 5'd6};
    assign wire4091 = {5'd12, 5'd6};
    assign wire4092 = {5'd12, 5'd6};
    assign wire4093 = {5'd12, 5'd6};
    assign wire4094 = {5'd12, 5'd6};
    assign wire4095 = {5'd12, 5'd6};
    wire [40959:0] data_concat;
    assign data_concat = {wire4095, wire4094, wire4093, wire4092, wire4091, wire4090, wire4089, wire4088, wire4087, wire4086, wire4085, wire4084, wire4083, wire4082, wire4081, wire4080, wire4079, wire4078, wire4077, wire4076, wire4075, wire4074, wire4073, wire4072, wire4071, wire4070, wire4069, wire4068, wire4067, wire4066, wire4065, wire4064, wire4063, wire4062, wire4061, wire4060, wire4059, wire4058, wire4057, wire4056, wire4055, wire4054, wire4053, wire4052, wire4051, wire4050, wire4049, wire4048, wire4047, wire4046, wire4045, wire4044, wire4043, wire4042, wire4041, wire4040, wire4039, wire4038, wire4037, wire4036, wire4035, wire4034, wire4033, wire4032, wire4031, wire4030, wire4029, wire4028, wire4027, wire4026, wire4025, wire4024, wire4023, wire4022, wire4021, wire4020, wire4019, wire4018, wire4017, wire4016, wire4015, wire4014, wire4013, wire4012, wire4011, wire4010, wire4009, wire4008, wire4007, wire4006, wire4005, wire4004, wire4003, wire4002, wire4001, wire4000, wire3999, wire3998, wire3997, wire3996, wire3995, wire3994, wire3993, wire3992, wire3991, wire3990, wire3989, wire3988, wire3987, wire3986, wire3985, wire3984, wire3983, wire3982, wire3981, wire3980, wire3979, wire3978, wire3977, wire3976, wire3975, wire3974, wire3973, wire3972, wire3971, wire3970, wire3969, wire3968, wire3967, wire3966, wire3965, wire3964, wire3963, wire3962, wire3961, wire3960, wire3959, wire3958, wire3957, wire3956, wire3955, wire3954, wire3953, wire3952, wire3951, wire3950, wire3949, wire3948, wire3947, wire3946, wire3945, wire3944, wire3943, wire3942, wire3941, wire3940, wire3939, wire3938, wire3937, wire3936, wire3935, wire3934, wire3933, wire3932, wire3931, wire3930, wire3929, wire3928, wire3927, wire3926, wire3925, wire3924, wire3923, wire3922, wire3921, wire3920, wire3919, wire3918, wire3917, wire3916, wire3915, wire3914, wire3913, wire3912, wire3911, wire3910, wire3909, wire3908, wire3907, wire3906, wire3905, wire3904, wire3903, wire3902, wire3901, wire3900, wire3899, wire3898, wire3897, wire3896, wire3895, wire3894, wire3893, wire3892, wire3891, wire3890, wire3889, wire3888, wire3887, wire3886, wire3885, wire3884, wire3883, wire3882, wire3881, wire3880, wire3879, wire3878, wire3877, wire3876, wire3875, wire3874, wire3873, wire3872, wire3871, wire3870, wire3869, wire3868, wire3867, wire3866, wire3865, wire3864, wire3863, wire3862, wire3861, wire3860, wire3859, wire3858, wire3857, wire3856, wire3855, wire3854, wire3853, wire3852, wire3851, wire3850, wire3849, wire3848, wire3847, wire3846, wire3845, wire3844, wire3843, wire3842, wire3841, wire3840, wire3839, wire3838, wire3837, wire3836, wire3835, wire3834, wire3833, wire3832, wire3831, wire3830, wire3829, wire3828, wire3827, wire3826, wire3825, wire3824, wire3823, wire3822, wire3821, wire3820, wire3819, wire3818, wire3817, wire3816, wire3815, wire3814, wire3813, wire3812, wire3811, wire3810, wire3809, wire3808, wire3807, wire3806, wire3805, wire3804, wire3803, wire3802, wire3801, wire3800, wire3799, wire3798, wire3797, wire3796, wire3795, wire3794, wire3793, wire3792, wire3791, wire3790, wire3789, wire3788, wire3787, wire3786, wire3785, wire3784, wire3783, wire3782, wire3781, wire3780, wire3779, wire3778, wire3777, wire3776, wire3775, wire3774, wire3773, wire3772, wire3771, wire3770, wire3769, wire3768, wire3767, wire3766, wire3765, wire3764, wire3763, wire3762, wire3761, wire3760, wire3759, wire3758, wire3757, wire3756, wire3755, wire3754, wire3753, wire3752, wire3751, wire3750, wire3749, wire3748, wire3747, wire3746, wire3745, wire3744, wire3743, wire3742, wire3741, wire3740, wire3739, wire3738, wire3737, wire3736, wire3735, wire3734, wire3733, wire3732, wire3731, wire3730, wire3729, wire3728, wire3727, wire3726, wire3725, wire3724, wire3723, wire3722, wire3721, wire3720, wire3719, wire3718, wire3717, wire3716, wire3715, wire3714, wire3713, wire3712, wire3711, wire3710, wire3709, wire3708, wire3707, wire3706, wire3705, wire3704, wire3703, wire3702, wire3701, wire3700, wire3699, wire3698, wire3697, wire3696, wire3695, wire3694, wire3693, wire3692, wire3691, wire3690, wire3689, wire3688, wire3687, wire3686, wire3685, wire3684, wire3683, wire3682, wire3681, wire3680, wire3679, wire3678, wire3677, wire3676, wire3675, wire3674, wire3673, wire3672, wire3671, wire3670, wire3669, wire3668, wire3667, wire3666, wire3665, wire3664, wire3663, wire3662, wire3661, wire3660, wire3659, wire3658, wire3657, wire3656, wire3655, wire3654, wire3653, wire3652, wire3651, wire3650, wire3649, wire3648, wire3647, wire3646, wire3645, wire3644, wire3643, wire3642, wire3641, wire3640, wire3639, wire3638, wire3637, wire3636, wire3635, wire3634, wire3633, wire3632, wire3631, wire3630, wire3629, wire3628, wire3627, wire3626, wire3625, wire3624, wire3623, wire3622, wire3621, wire3620, wire3619, wire3618, wire3617, wire3616, wire3615, wire3614, wire3613, wire3612, wire3611, wire3610, wire3609, wire3608, wire3607, wire3606, wire3605, wire3604, wire3603, wire3602, wire3601, wire3600, wire3599, wire3598, wire3597, wire3596, wire3595, wire3594, wire3593, wire3592, wire3591, wire3590, wire3589, wire3588, wire3587, wire3586, wire3585, wire3584, wire3583, wire3582, wire3581, wire3580, wire3579, wire3578, wire3577, wire3576, wire3575, wire3574, wire3573, wire3572, wire3571, wire3570, wire3569, wire3568, wire3567, wire3566, wire3565, wire3564, wire3563, wire3562, wire3561, wire3560, wire3559, wire3558, wire3557, wire3556, wire3555, wire3554, wire3553, wire3552, wire3551, wire3550, wire3549, wire3548, wire3547, wire3546, wire3545, wire3544, wire3543, wire3542, wire3541, wire3540, wire3539, wire3538, wire3537, wire3536, wire3535, wire3534, wire3533, wire3532, wire3531, wire3530, wire3529, wire3528, wire3527, wire3526, wire3525, wire3524, wire3523, wire3522, wire3521, wire3520, wire3519, wire3518, wire3517, wire3516, wire3515, wire3514, wire3513, wire3512, wire3511, wire3510, wire3509, wire3508, wire3507, wire3506, wire3505, wire3504, wire3503, wire3502, wire3501, wire3500, wire3499, wire3498, wire3497, wire3496, wire3495, wire3494, wire3493, wire3492, wire3491, wire3490, wire3489, wire3488, wire3487, wire3486, wire3485, wire3484, wire3483, wire3482, wire3481, wire3480, wire3479, wire3478, wire3477, wire3476, wire3475, wire3474, wire3473, wire3472, wire3471, wire3470, wire3469, wire3468, wire3467, wire3466, wire3465, wire3464, wire3463, wire3462, wire3461, wire3460, wire3459, wire3458, wire3457, wire3456, wire3455, wire3454, wire3453, wire3452, wire3451, wire3450, wire3449, wire3448, wire3447, wire3446, wire3445, wire3444, wire3443, wire3442, wire3441, wire3440, wire3439, wire3438, wire3437, wire3436, wire3435, wire3434, wire3433, wire3432, wire3431, wire3430, wire3429, wire3428, wire3427, wire3426, wire3425, wire3424, wire3423, wire3422, wire3421, wire3420, wire3419, wire3418, wire3417, wire3416, wire3415, wire3414, wire3413, wire3412, wire3411, wire3410, wire3409, wire3408, wire3407, wire3406, wire3405, wire3404, wire3403, wire3402, wire3401, wire3400, wire3399, wire3398, wire3397, wire3396, wire3395, wire3394, wire3393, wire3392, wire3391, wire3390, wire3389, wire3388, wire3387, wire3386, wire3385, wire3384, wire3383, wire3382, wire3381, wire3380, wire3379, wire3378, wire3377, wire3376, wire3375, wire3374, wire3373, wire3372, wire3371, wire3370, wire3369, wire3368, wire3367, wire3366, wire3365, wire3364, wire3363, wire3362, wire3361, wire3360, wire3359, wire3358, wire3357, wire3356, wire3355, wire3354, wire3353, wire3352, wire3351, wire3350, wire3349, wire3348, wire3347, wire3346, wire3345, wire3344, wire3343, wire3342, wire3341, wire3340, wire3339, wire3338, wire3337, wire3336, wire3335, wire3334, wire3333, wire3332, wire3331, wire3330, wire3329, wire3328, wire3327, wire3326, wire3325, wire3324, wire3323, wire3322, wire3321, wire3320, wire3319, wire3318, wire3317, wire3316, wire3315, wire3314, wire3313, wire3312, wire3311, wire3310, wire3309, wire3308, wire3307, wire3306, wire3305, wire3304, wire3303, wire3302, wire3301, wire3300, wire3299, wire3298, wire3297, wire3296, wire3295, wire3294, wire3293, wire3292, wire3291, wire3290, wire3289, wire3288, wire3287, wire3286, wire3285, wire3284, wire3283, wire3282, wire3281, wire3280, wire3279, wire3278, wire3277, wire3276, wire3275, wire3274, wire3273, wire3272, wire3271, wire3270, wire3269, wire3268, wire3267, wire3266, wire3265, wire3264, wire3263, wire3262, wire3261, wire3260, wire3259, wire3258, wire3257, wire3256, wire3255, wire3254, wire3253, wire3252, wire3251, wire3250, wire3249, wire3248, wire3247, wire3246, wire3245, wire3244, wire3243, wire3242, wire3241, wire3240, wire3239, wire3238, wire3237, wire3236, wire3235, wire3234, wire3233, wire3232, wire3231, wire3230, wire3229, wire3228, wire3227, wire3226, wire3225, wire3224, wire3223, wire3222, wire3221, wire3220, wire3219, wire3218, wire3217, wire3216, wire3215, wire3214, wire3213, wire3212, wire3211, wire3210, wire3209, wire3208, wire3207, wire3206, wire3205, wire3204, wire3203, wire3202, wire3201, wire3200, wire3199, wire3198, wire3197, wire3196, wire3195, wire3194, wire3193, wire3192, wire3191, wire3190, wire3189, wire3188, wire3187, wire3186, wire3185, wire3184, wire3183, wire3182, wire3181, wire3180, wire3179, wire3178, wire3177, wire3176, wire3175, wire3174, wire3173, wire3172, wire3171, wire3170, wire3169, wire3168, wire3167, wire3166, wire3165, wire3164, wire3163, wire3162, wire3161, wire3160, wire3159, wire3158, wire3157, wire3156, wire3155, wire3154, wire3153, wire3152, wire3151, wire3150, wire3149, wire3148, wire3147, wire3146, wire3145, wire3144, wire3143, wire3142, wire3141, wire3140, wire3139, wire3138, wire3137, wire3136, wire3135, wire3134, wire3133, wire3132, wire3131, wire3130, wire3129, wire3128, wire3127, wire3126, wire3125, wire3124, wire3123, wire3122, wire3121, wire3120, wire3119, wire3118, wire3117, wire3116, wire3115, wire3114, wire3113, wire3112, wire3111, wire3110, wire3109, wire3108, wire3107, wire3106, wire3105, wire3104, wire3103, wire3102, wire3101, wire3100, wire3099, wire3098, wire3097, wire3096, wire3095, wire3094, wire3093, wire3092, wire3091, wire3090, wire3089, wire3088, wire3087, wire3086, wire3085, wire3084, wire3083, wire3082, wire3081, wire3080, wire3079, wire3078, wire3077, wire3076, wire3075, wire3074, wire3073, wire3072, wire3071, wire3070, wire3069, wire3068, wire3067, wire3066, wire3065, wire3064, wire3063, wire3062, wire3061, wire3060, wire3059, wire3058, wire3057, wire3056, wire3055, wire3054, wire3053, wire3052, wire3051, wire3050, wire3049, wire3048, wire3047, wire3046, wire3045, wire3044, wire3043, wire3042, wire3041, wire3040, wire3039, wire3038, wire3037, wire3036, wire3035, wire3034, wire3033, wire3032, wire3031, wire3030, wire3029, wire3028, wire3027, wire3026, wire3025, wire3024, wire3023, wire3022, wire3021, wire3020, wire3019, wire3018, wire3017, wire3016, wire3015, wire3014, wire3013, wire3012, wire3011, wire3010, wire3009, wire3008, wire3007, wire3006, wire3005, wire3004, wire3003, wire3002, wire3001, wire3000, wire2999, wire2998, wire2997, wire2996, wire2995, wire2994, wire2993, wire2992, wire2991, wire2990, wire2989, wire2988, wire2987, wire2986, wire2985, wire2984, wire2983, wire2982, wire2981, wire2980, wire2979, wire2978, wire2977, wire2976, wire2975, wire2974, wire2973, wire2972, wire2971, wire2970, wire2969, wire2968, wire2967, wire2966, wire2965, wire2964, wire2963, wire2962, wire2961, wire2960, wire2959, wire2958, wire2957, wire2956, wire2955, wire2954, wire2953, wire2952, wire2951, wire2950, wire2949, wire2948, wire2947, wire2946, wire2945, wire2944, wire2943, wire2942, wire2941, wire2940, wire2939, wire2938, wire2937, wire2936, wire2935, wire2934, wire2933, wire2932, wire2931, wire2930, wire2929, wire2928, wire2927, wire2926, wire2925, wire2924, wire2923, wire2922, wire2921, wire2920, wire2919, wire2918, wire2917, wire2916, wire2915, wire2914, wire2913, wire2912, wire2911, wire2910, wire2909, wire2908, wire2907, wire2906, wire2905, wire2904, wire2903, wire2902, wire2901, wire2900, wire2899, wire2898, wire2897, wire2896, wire2895, wire2894, wire2893, wire2892, wire2891, wire2890, wire2889, wire2888, wire2887, wire2886, wire2885, wire2884, wire2883, wire2882, wire2881, wire2880, wire2879, wire2878, wire2877, wire2876, wire2875, wire2874, wire2873, wire2872, wire2871, wire2870, wire2869, wire2868, wire2867, wire2866, wire2865, wire2864, wire2863, wire2862, wire2861, wire2860, wire2859, wire2858, wire2857, wire2856, wire2855, wire2854, wire2853, wire2852, wire2851, wire2850, wire2849, wire2848, wire2847, wire2846, wire2845, wire2844, wire2843, wire2842, wire2841, wire2840, wire2839, wire2838, wire2837, wire2836, wire2835, wire2834, wire2833, wire2832, wire2831, wire2830, wire2829, wire2828, wire2827, wire2826, wire2825, wire2824, wire2823, wire2822, wire2821, wire2820, wire2819, wire2818, wire2817, wire2816, wire2815, wire2814, wire2813, wire2812, wire2811, wire2810, wire2809, wire2808, wire2807, wire2806, wire2805, wire2804, wire2803, wire2802, wire2801, wire2800, wire2799, wire2798, wire2797, wire2796, wire2795, wire2794, wire2793, wire2792, wire2791, wire2790, wire2789, wire2788, wire2787, wire2786, wire2785, wire2784, wire2783, wire2782, wire2781, wire2780, wire2779, wire2778, wire2777, wire2776, wire2775, wire2774, wire2773, wire2772, wire2771, wire2770, wire2769, wire2768, wire2767, wire2766, wire2765, wire2764, wire2763, wire2762, wire2761, wire2760, wire2759, wire2758, wire2757, wire2756, wire2755, wire2754, wire2753, wire2752, wire2751, wire2750, wire2749, wire2748, wire2747, wire2746, wire2745, wire2744, wire2743, wire2742, wire2741, wire2740, wire2739, wire2738, wire2737, wire2736, wire2735, wire2734, wire2733, wire2732, wire2731, wire2730, wire2729, wire2728, wire2727, wire2726, wire2725, wire2724, wire2723, wire2722, wire2721, wire2720, wire2719, wire2718, wire2717, wire2716, wire2715, wire2714, wire2713, wire2712, wire2711, wire2710, wire2709, wire2708, wire2707, wire2706, wire2705, wire2704, wire2703, wire2702, wire2701, wire2700, wire2699, wire2698, wire2697, wire2696, wire2695, wire2694, wire2693, wire2692, wire2691, wire2690, wire2689, wire2688, wire2687, wire2686, wire2685, wire2684, wire2683, wire2682, wire2681, wire2680, wire2679, wire2678, wire2677, wire2676, wire2675, wire2674, wire2673, wire2672, wire2671, wire2670, wire2669, wire2668, wire2667, wire2666, wire2665, wire2664, wire2663, wire2662, wire2661, wire2660, wire2659, wire2658, wire2657, wire2656, wire2655, wire2654, wire2653, wire2652, wire2651, wire2650, wire2649, wire2648, wire2647, wire2646, wire2645, wire2644, wire2643, wire2642, wire2641, wire2640, wire2639, wire2638, wire2637, wire2636, wire2635, wire2634, wire2633, wire2632, wire2631, wire2630, wire2629, wire2628, wire2627, wire2626, wire2625, wire2624, wire2623, wire2622, wire2621, wire2620, wire2619, wire2618, wire2617, wire2616, wire2615, wire2614, wire2613, wire2612, wire2611, wire2610, wire2609, wire2608, wire2607, wire2606, wire2605, wire2604, wire2603, wire2602, wire2601, wire2600, wire2599, wire2598, wire2597, wire2596, wire2595, wire2594, wire2593, wire2592, wire2591, wire2590, wire2589, wire2588, wire2587, wire2586, wire2585, wire2584, wire2583, wire2582, wire2581, wire2580, wire2579, wire2578, wire2577, wire2576, wire2575, wire2574, wire2573, wire2572, wire2571, wire2570, wire2569, wire2568, wire2567, wire2566, wire2565, wire2564, wire2563, wire2562, wire2561, wire2560, wire2559, wire2558, wire2557, wire2556, wire2555, wire2554, wire2553, wire2552, wire2551, wire2550, wire2549, wire2548, wire2547, wire2546, wire2545, wire2544, wire2543, wire2542, wire2541, wire2540, wire2539, wire2538, wire2537, wire2536, wire2535, wire2534, wire2533, wire2532, wire2531, wire2530, wire2529, wire2528, wire2527, wire2526, wire2525, wire2524, wire2523, wire2522, wire2521, wire2520, wire2519, wire2518, wire2517, wire2516, wire2515, wire2514, wire2513, wire2512, wire2511, wire2510, wire2509, wire2508, wire2507, wire2506, wire2505, wire2504, wire2503, wire2502, wire2501, wire2500, wire2499, wire2498, wire2497, wire2496, wire2495, wire2494, wire2493, wire2492, wire2491, wire2490, wire2489, wire2488, wire2487, wire2486, wire2485, wire2484, wire2483, wire2482, wire2481, wire2480, wire2479, wire2478, wire2477, wire2476, wire2475, wire2474, wire2473, wire2472, wire2471, wire2470, wire2469, wire2468, wire2467, wire2466, wire2465, wire2464, wire2463, wire2462, wire2461, wire2460, wire2459, wire2458, wire2457, wire2456, wire2455, wire2454, wire2453, wire2452, wire2451, wire2450, wire2449, wire2448, wire2447, wire2446, wire2445, wire2444, wire2443, wire2442, wire2441, wire2440, wire2439, wire2438, wire2437, wire2436, wire2435, wire2434, wire2433, wire2432, wire2431, wire2430, wire2429, wire2428, wire2427, wire2426, wire2425, wire2424, wire2423, wire2422, wire2421, wire2420, wire2419, wire2418, wire2417, wire2416, wire2415, wire2414, wire2413, wire2412, wire2411, wire2410, wire2409, wire2408, wire2407, wire2406, wire2405, wire2404, wire2403, wire2402, wire2401, wire2400, wire2399, wire2398, wire2397, wire2396, wire2395, wire2394, wire2393, wire2392, wire2391, wire2390, wire2389, wire2388, wire2387, wire2386, wire2385, wire2384, wire2383, wire2382, wire2381, wire2380, wire2379, wire2378, wire2377, wire2376, wire2375, wire2374, wire2373, wire2372, wire2371, wire2370, wire2369, wire2368, wire2367, wire2366, wire2365, wire2364, wire2363, wire2362, wire2361, wire2360, wire2359, wire2358, wire2357, wire2356, wire2355, wire2354, wire2353, wire2352, wire2351, wire2350, wire2349, wire2348, wire2347, wire2346, wire2345, wire2344, wire2343, wire2342, wire2341, wire2340, wire2339, wire2338, wire2337, wire2336, wire2335, wire2334, wire2333, wire2332, wire2331, wire2330, wire2329, wire2328, wire2327, wire2326, wire2325, wire2324, wire2323, wire2322, wire2321, wire2320, wire2319, wire2318, wire2317, wire2316, wire2315, wire2314, wire2313, wire2312, wire2311, wire2310, wire2309, wire2308, wire2307, wire2306, wire2305, wire2304, wire2303, wire2302, wire2301, wire2300, wire2299, wire2298, wire2297, wire2296, wire2295, wire2294, wire2293, wire2292, wire2291, wire2290, wire2289, wire2288, wire2287, wire2286, wire2285, wire2284, wire2283, wire2282, wire2281, wire2280, wire2279, wire2278, wire2277, wire2276, wire2275, wire2274, wire2273, wire2272, wire2271, wire2270, wire2269, wire2268, wire2267, wire2266, wire2265, wire2264, wire2263, wire2262, wire2261, wire2260, wire2259, wire2258, wire2257, wire2256, wire2255, wire2254, wire2253, wire2252, wire2251, wire2250, wire2249, wire2248, wire2247, wire2246, wire2245, wire2244, wire2243, wire2242, wire2241, wire2240, wire2239, wire2238, wire2237, wire2236, wire2235, wire2234, wire2233, wire2232, wire2231, wire2230, wire2229, wire2228, wire2227, wire2226, wire2225, wire2224, wire2223, wire2222, wire2221, wire2220, wire2219, wire2218, wire2217, wire2216, wire2215, wire2214, wire2213, wire2212, wire2211, wire2210, wire2209, wire2208, wire2207, wire2206, wire2205, wire2204, wire2203, wire2202, wire2201, wire2200, wire2199, wire2198, wire2197, wire2196, wire2195, wire2194, wire2193, wire2192, wire2191, wire2190, wire2189, wire2188, wire2187, wire2186, wire2185, wire2184, wire2183, wire2182, wire2181, wire2180, wire2179, wire2178, wire2177, wire2176, wire2175, wire2174, wire2173, wire2172, wire2171, wire2170, wire2169, wire2168, wire2167, wire2166, wire2165, wire2164, wire2163, wire2162, wire2161, wire2160, wire2159, wire2158, wire2157, wire2156, wire2155, wire2154, wire2153, wire2152, wire2151, wire2150, wire2149, wire2148, wire2147, wire2146, wire2145, wire2144, wire2143, wire2142, wire2141, wire2140, wire2139, wire2138, wire2137, wire2136, wire2135, wire2134, wire2133, wire2132, wire2131, wire2130, wire2129, wire2128, wire2127, wire2126, wire2125, wire2124, wire2123, wire2122, wire2121, wire2120, wire2119, wire2118, wire2117, wire2116, wire2115, wire2114, wire2113, wire2112, wire2111, wire2110, wire2109, wire2108, wire2107, wire2106, wire2105, wire2104, wire2103, wire2102, wire2101, wire2100, wire2099, wire2098, wire2097, wire2096, wire2095, wire2094, wire2093, wire2092, wire2091, wire2090, wire2089, wire2088, wire2087, wire2086, wire2085, wire2084, wire2083, wire2082, wire2081, wire2080, wire2079, wire2078, wire2077, wire2076, wire2075, wire2074, wire2073, wire2072, wire2071, wire2070, wire2069, wire2068, wire2067, wire2066, wire2065, wire2064, wire2063, wire2062, wire2061, wire2060, wire2059, wire2058, wire2057, wire2056, wire2055, wire2054, wire2053, wire2052, wire2051, wire2050, wire2049, wire2048, wire2047, wire2046, wire2045, wire2044, wire2043, wire2042, wire2041, wire2040, wire2039, wire2038, wire2037, wire2036, wire2035, wire2034, wire2033, wire2032, wire2031, wire2030, wire2029, wire2028, wire2027, wire2026, wire2025, wire2024, wire2023, wire2022, wire2021, wire2020, wire2019, wire2018, wire2017, wire2016, wire2015, wire2014, wire2013, wire2012, wire2011, wire2010, wire2009, wire2008, wire2007, wire2006, wire2005, wire2004, wire2003, wire2002, wire2001, wire2000, wire1999, wire1998, wire1997, wire1996, wire1995, wire1994, wire1993, wire1992, wire1991, wire1990, wire1989, wire1988, wire1987, wire1986, wire1985, wire1984, wire1983, wire1982, wire1981, wire1980, wire1979, wire1978, wire1977, wire1976, wire1975, wire1974, wire1973, wire1972, wire1971, wire1970, wire1969, wire1968, wire1967, wire1966, wire1965, wire1964, wire1963, wire1962, wire1961, wire1960, wire1959, wire1958, wire1957, wire1956, wire1955, wire1954, wire1953, wire1952, wire1951, wire1950, wire1949, wire1948, wire1947, wire1946, wire1945, wire1944, wire1943, wire1942, wire1941, wire1940, wire1939, wire1938, wire1937, wire1936, wire1935, wire1934, wire1933, wire1932, wire1931, wire1930, wire1929, wire1928, wire1927, wire1926, wire1925, wire1924, wire1923, wire1922, wire1921, wire1920, wire1919, wire1918, wire1917, wire1916, wire1915, wire1914, wire1913, wire1912, wire1911, wire1910, wire1909, wire1908, wire1907, wire1906, wire1905, wire1904, wire1903, wire1902, wire1901, wire1900, wire1899, wire1898, wire1897, wire1896, wire1895, wire1894, wire1893, wire1892, wire1891, wire1890, wire1889, wire1888, wire1887, wire1886, wire1885, wire1884, wire1883, wire1882, wire1881, wire1880, wire1879, wire1878, wire1877, wire1876, wire1875, wire1874, wire1873, wire1872, wire1871, wire1870, wire1869, wire1868, wire1867, wire1866, wire1865, wire1864, wire1863, wire1862, wire1861, wire1860, wire1859, wire1858, wire1857, wire1856, wire1855, wire1854, wire1853, wire1852, wire1851, wire1850, wire1849, wire1848, wire1847, wire1846, wire1845, wire1844, wire1843, wire1842, wire1841, wire1840, wire1839, wire1838, wire1837, wire1836, wire1835, wire1834, wire1833, wire1832, wire1831, wire1830, wire1829, wire1828, wire1827, wire1826, wire1825, wire1824, wire1823, wire1822, wire1821, wire1820, wire1819, wire1818, wire1817, wire1816, wire1815, wire1814, wire1813, wire1812, wire1811, wire1810, wire1809, wire1808, wire1807, wire1806, wire1805, wire1804, wire1803, wire1802, wire1801, wire1800, wire1799, wire1798, wire1797, wire1796, wire1795, wire1794, wire1793, wire1792, wire1791, wire1790, wire1789, wire1788, wire1787, wire1786, wire1785, wire1784, wire1783, wire1782, wire1781, wire1780, wire1779, wire1778, wire1777, wire1776, wire1775, wire1774, wire1773, wire1772, wire1771, wire1770, wire1769, wire1768, wire1767, wire1766, wire1765, wire1764, wire1763, wire1762, wire1761, wire1760, wire1759, wire1758, wire1757, wire1756, wire1755, wire1754, wire1753, wire1752, wire1751, wire1750, wire1749, wire1748, wire1747, wire1746, wire1745, wire1744, wire1743, wire1742, wire1741, wire1740, wire1739, wire1738, wire1737, wire1736, wire1735, wire1734, wire1733, wire1732, wire1731, wire1730, wire1729, wire1728, wire1727, wire1726, wire1725, wire1724, wire1723, wire1722, wire1721, wire1720, wire1719, wire1718, wire1717, wire1716, wire1715, wire1714, wire1713, wire1712, wire1711, wire1710, wire1709, wire1708, wire1707, wire1706, wire1705, wire1704, wire1703, wire1702, wire1701, wire1700, wire1699, wire1698, wire1697, wire1696, wire1695, wire1694, wire1693, wire1692, wire1691, wire1690, wire1689, wire1688, wire1687, wire1686, wire1685, wire1684, wire1683, wire1682, wire1681, wire1680, wire1679, wire1678, wire1677, wire1676, wire1675, wire1674, wire1673, wire1672, wire1671, wire1670, wire1669, wire1668, wire1667, wire1666, wire1665, wire1664, wire1663, wire1662, wire1661, wire1660, wire1659, wire1658, wire1657, wire1656, wire1655, wire1654, wire1653, wire1652, wire1651, wire1650, wire1649, wire1648, wire1647, wire1646, wire1645, wire1644, wire1643, wire1642, wire1641, wire1640, wire1639, wire1638, wire1637, wire1636, wire1635, wire1634, wire1633, wire1632, wire1631, wire1630, wire1629, wire1628, wire1627, wire1626, wire1625, wire1624, wire1623, wire1622, wire1621, wire1620, wire1619, wire1618, wire1617, wire1616, wire1615, wire1614, wire1613, wire1612, wire1611, wire1610, wire1609, wire1608, wire1607, wire1606, wire1605, wire1604, wire1603, wire1602, wire1601, wire1600, wire1599, wire1598, wire1597, wire1596, wire1595, wire1594, wire1593, wire1592, wire1591, wire1590, wire1589, wire1588, wire1587, wire1586, wire1585, wire1584, wire1583, wire1582, wire1581, wire1580, wire1579, wire1578, wire1577, wire1576, wire1575, wire1574, wire1573, wire1572, wire1571, wire1570, wire1569, wire1568, wire1567, wire1566, wire1565, wire1564, wire1563, wire1562, wire1561, wire1560, wire1559, wire1558, wire1557, wire1556, wire1555, wire1554, wire1553, wire1552, wire1551, wire1550, wire1549, wire1548, wire1547, wire1546, wire1545, wire1544, wire1543, wire1542, wire1541, wire1540, wire1539, wire1538, wire1537, wire1536, wire1535, wire1534, wire1533, wire1532, wire1531, wire1530, wire1529, wire1528, wire1527, wire1526, wire1525, wire1524, wire1523, wire1522, wire1521, wire1520, wire1519, wire1518, wire1517, wire1516, wire1515, wire1514, wire1513, wire1512, wire1511, wire1510, wire1509, wire1508, wire1507, wire1506, wire1505, wire1504, wire1503, wire1502, wire1501, wire1500, wire1499, wire1498, wire1497, wire1496, wire1495, wire1494, wire1493, wire1492, wire1491, wire1490, wire1489, wire1488, wire1487, wire1486, wire1485, wire1484, wire1483, wire1482, wire1481, wire1480, wire1479, wire1478, wire1477, wire1476, wire1475, wire1474, wire1473, wire1472, wire1471, wire1470, wire1469, wire1468, wire1467, wire1466, wire1465, wire1464, wire1463, wire1462, wire1461, wire1460, wire1459, wire1458, wire1457, wire1456, wire1455, wire1454, wire1453, wire1452, wire1451, wire1450, wire1449, wire1448, wire1447, wire1446, wire1445, wire1444, wire1443, wire1442, wire1441, wire1440, wire1439, wire1438, wire1437, wire1436, wire1435, wire1434, wire1433, wire1432, wire1431, wire1430, wire1429, wire1428, wire1427, wire1426, wire1425, wire1424, wire1423, wire1422, wire1421, wire1420, wire1419, wire1418, wire1417, wire1416, wire1415, wire1414, wire1413, wire1412, wire1411, wire1410, wire1409, wire1408, wire1407, wire1406, wire1405, wire1404, wire1403, wire1402, wire1401, wire1400, wire1399, wire1398, wire1397, wire1396, wire1395, wire1394, wire1393, wire1392, wire1391, wire1390, wire1389, wire1388, wire1387, wire1386, wire1385, wire1384, wire1383, wire1382, wire1381, wire1380, wire1379, wire1378, wire1377, wire1376, wire1375, wire1374, wire1373, wire1372, wire1371, wire1370, wire1369, wire1368, wire1367, wire1366, wire1365, wire1364, wire1363, wire1362, wire1361, wire1360, wire1359, wire1358, wire1357, wire1356, wire1355, wire1354, wire1353, wire1352, wire1351, wire1350, wire1349, wire1348, wire1347, wire1346, wire1345, wire1344, wire1343, wire1342, wire1341, wire1340, wire1339, wire1338, wire1337, wire1336, wire1335, wire1334, wire1333, wire1332, wire1331, wire1330, wire1329, wire1328, wire1327, wire1326, wire1325, wire1324, wire1323, wire1322, wire1321, wire1320, wire1319, wire1318, wire1317, wire1316, wire1315, wire1314, wire1313, wire1312, wire1311, wire1310, wire1309, wire1308, wire1307, wire1306, wire1305, wire1304, wire1303, wire1302, wire1301, wire1300, wire1299, wire1298, wire1297, wire1296, wire1295, wire1294, wire1293, wire1292, wire1291, wire1290, wire1289, wire1288, wire1287, wire1286, wire1285, wire1284, wire1283, wire1282, wire1281, wire1280, wire1279, wire1278, wire1277, wire1276, wire1275, wire1274, wire1273, wire1272, wire1271, wire1270, wire1269, wire1268, wire1267, wire1266, wire1265, wire1264, wire1263, wire1262, wire1261, wire1260, wire1259, wire1258, wire1257, wire1256, wire1255, wire1254, wire1253, wire1252, wire1251, wire1250, wire1249, wire1248, wire1247, wire1246, wire1245, wire1244, wire1243, wire1242, wire1241, wire1240, wire1239, wire1238, wire1237, wire1236, wire1235, wire1234, wire1233, wire1232, wire1231, wire1230, wire1229, wire1228, wire1227, wire1226, wire1225, wire1224, wire1223, wire1222, wire1221, wire1220, wire1219, wire1218, wire1217, wire1216, wire1215, wire1214, wire1213, wire1212, wire1211, wire1210, wire1209, wire1208, wire1207, wire1206, wire1205, wire1204, wire1203, wire1202, wire1201, wire1200, wire1199, wire1198, wire1197, wire1196, wire1195, wire1194, wire1193, wire1192, wire1191, wire1190, wire1189, wire1188, wire1187, wire1186, wire1185, wire1184, wire1183, wire1182, wire1181, wire1180, wire1179, wire1178, wire1177, wire1176, wire1175, wire1174, wire1173, wire1172, wire1171, wire1170, wire1169, wire1168, wire1167, wire1166, wire1165, wire1164, wire1163, wire1162, wire1161, wire1160, wire1159, wire1158, wire1157, wire1156, wire1155, wire1154, wire1153, wire1152, wire1151, wire1150, wire1149, wire1148, wire1147, wire1146, wire1145, wire1144, wire1143, wire1142, wire1141, wire1140, wire1139, wire1138, wire1137, wire1136, wire1135, wire1134, wire1133, wire1132, wire1131, wire1130, wire1129, wire1128, wire1127, wire1126, wire1125, wire1124, wire1123, wire1122, wire1121, wire1120, wire1119, wire1118, wire1117, wire1116, wire1115, wire1114, wire1113, wire1112, wire1111, wire1110, wire1109, wire1108, wire1107, wire1106, wire1105, wire1104, wire1103, wire1102, wire1101, wire1100, wire1099, wire1098, wire1097, wire1096, wire1095, wire1094, wire1093, wire1092, wire1091, wire1090, wire1089, wire1088, wire1087, wire1086, wire1085, wire1084, wire1083, wire1082, wire1081, wire1080, wire1079, wire1078, wire1077, wire1076, wire1075, wire1074, wire1073, wire1072, wire1071, wire1070, wire1069, wire1068, wire1067, wire1066, wire1065, wire1064, wire1063, wire1062, wire1061, wire1060, wire1059, wire1058, wire1057, wire1056, wire1055, wire1054, wire1053, wire1052, wire1051, wire1050, wire1049, wire1048, wire1047, wire1046, wire1045, wire1044, wire1043, wire1042, wire1041, wire1040, wire1039, wire1038, wire1037, wire1036, wire1035, wire1034, wire1033, wire1032, wire1031, wire1030, wire1029, wire1028, wire1027, wire1026, wire1025, wire1024, wire1023, wire1022, wire1021, wire1020, wire1019, wire1018, wire1017, wire1016, wire1015, wire1014, wire1013, wire1012, wire1011, wire1010, wire1009, wire1008, wire1007, wire1006, wire1005, wire1004, wire1003, wire1002, wire1001, wire1000, wire999, wire998, wire997, wire996, wire995, wire994, wire993, wire992, wire991, wire990, wire989, wire988, wire987, wire986, wire985, wire984, wire983, wire982, wire981, wire980, wire979, wire978, wire977, wire976, wire975, wire974, wire973, wire972, wire971, wire970, wire969, wire968, wire967, wire966, wire965, wire964, wire963, wire962, wire961, wire960, wire959, wire958, wire957, wire956, wire955, wire954, wire953, wire952, wire951, wire950, wire949, wire948, wire947, wire946, wire945, wire944, wire943, wire942, wire941, wire940, wire939, wire938, wire937, wire936, wire935, wire934, wire933, wire932, wire931, wire930, wire929, wire928, wire927, wire926, wire925, wire924, wire923, wire922, wire921, wire920, wire919, wire918, wire917, wire916, wire915, wire914, wire913, wire912, wire911, wire910, wire909, wire908, wire907, wire906, wire905, wire904, wire903, wire902, wire901, wire900, wire899, wire898, wire897, wire896, wire895, wire894, wire893, wire892, wire891, wire890, wire889, wire888, wire887, wire886, wire885, wire884, wire883, wire882, wire881, wire880, wire879, wire878, wire877, wire876, wire875, wire874, wire873, wire872, wire871, wire870, wire869, wire868, wire867, wire866, wire865, wire864, wire863, wire862, wire861, wire860, wire859, wire858, wire857, wire856, wire855, wire854, wire853, wire852, wire851, wire850, wire849, wire848, wire847, wire846, wire845, wire844, wire843, wire842, wire841, wire840, wire839, wire838, wire837, wire836, wire835, wire834, wire833, wire832, wire831, wire830, wire829, wire828, wire827, wire826, wire825, wire824, wire823, wire822, wire821, wire820, wire819, wire818, wire817, wire816, wire815, wire814, wire813, wire812, wire811, wire810, wire809, wire808, wire807, wire806, wire805, wire804, wire803, wire802, wire801, wire800, wire799, wire798, wire797, wire796, wire795, wire794, wire793, wire792, wire791, wire790, wire789, wire788, wire787, wire786, wire785, wire784, wire783, wire782, wire781, wire780, wire779, wire778, wire777, wire776, wire775, wire774, wire773, wire772, wire771, wire770, wire769, wire768, wire767, wire766, wire765, wire764, wire763, wire762, wire761, wire760, wire759, wire758, wire757, wire756, wire755, wire754, wire753, wire752, wire751, wire750, wire749, wire748, wire747, wire746, wire745, wire744, wire743, wire742, wire741, wire740, wire739, wire738, wire737, wire736, wire735, wire734, wire733, wire732, wire731, wire730, wire729, wire728, wire727, wire726, wire725, wire724, wire723, wire722, wire721, wire720, wire719, wire718, wire717, wire716, wire715, wire714, wire713, wire712, wire711, wire710, wire709, wire708, wire707, wire706, wire705, wire704, wire703, wire702, wire701, wire700, wire699, wire698, wire697, wire696, wire695, wire694, wire693, wire692, wire691, wire690, wire689, wire688, wire687, wire686, wire685, wire684, wire683, wire682, wire681, wire680, wire679, wire678, wire677, wire676, wire675, wire674, wire673, wire672, wire671, wire670, wire669, wire668, wire667, wire666, wire665, wire664, wire663, wire662, wire661, wire660, wire659, wire658, wire657, wire656, wire655, wire654, wire653, wire652, wire651, wire650, wire649, wire648, wire647, wire646, wire645, wire644, wire643, wire642, wire641, wire640, wire639, wire638, wire637, wire636, wire635, wire634, wire633, wire632, wire631, wire630, wire629, wire628, wire627, wire626, wire625, wire624, wire623, wire622, wire621, wire620, wire619, wire618, wire617, wire616, wire615, wire614, wire613, wire612, wire611, wire610, wire609, wire608, wire607, wire606, wire605, wire604, wire603, wire602, wire601, wire600, wire599, wire598, wire597, wire596, wire595, wire594, wire593, wire592, wire591, wire590, wire589, wire588, wire587, wire586, wire585, wire584, wire583, wire582, wire581, wire580, wire579, wire578, wire577, wire576, wire575, wire574, wire573, wire572, wire571, wire570, wire569, wire568, wire567, wire566, wire565, wire564, wire563, wire562, wire561, wire560, wire559, wire558, wire557, wire556, wire555, wire554, wire553, wire552, wire551, wire550, wire549, wire548, wire547, wire546, wire545, wire544, wire543, wire542, wire541, wire540, wire539, wire538, wire537, wire536, wire535, wire534, wire533, wire532, wire531, wire530, wire529, wire528, wire527, wire526, wire525, wire524, wire523, wire522, wire521, wire520, wire519, wire518, wire517, wire516, wire515, wire514, wire513, wire512, wire511, wire510, wire509, wire508, wire507, wire506, wire505, wire504, wire503, wire502, wire501, wire500, wire499, wire498, wire497, wire496, wire495, wire494, wire493, wire492, wire491, wire490, wire489, wire488, wire487, wire486, wire485, wire484, wire483, wire482, wire481, wire480, wire479, wire478, wire477, wire476, wire475, wire474, wire473, wire472, wire471, wire470, wire469, wire468, wire467, wire466, wire465, wire464, wire463, wire462, wire461, wire460, wire459, wire458, wire457, wire456, wire455, wire454, wire453, wire452, wire451, wire450, wire449, wire448, wire447, wire446, wire445, wire444, wire443, wire442, wire441, wire440, wire439, wire438, wire437, wire436, wire435, wire434, wire433, wire432, wire431, wire430, wire429, wire428, wire427, wire426, wire425, wire424, wire423, wire422, wire421, wire420, wire419, wire418, wire417, wire416, wire415, wire414, wire413, wire412, wire411, wire410, wire409, wire408, wire407, wire406, wire405, wire404, wire403, wire402, wire401, wire400, wire399, wire398, wire397, wire396, wire395, wire394, wire393, wire392, wire391, wire390, wire389, wire388, wire387, wire386, wire385, wire384, wire383, wire382, wire381, wire380, wire379, wire378, wire377, wire376, wire375, wire374, wire373, wire372, wire371, wire370, wire369, wire368, wire367, wire366, wire365, wire364, wire363, wire362, wire361, wire360, wire359, wire358, wire357, wire356, wire355, wire354, wire353, wire352, wire351, wire350, wire349, wire348, wire347, wire346, wire345, wire344, wire343, wire342, wire341, wire340, wire339, wire338, wire337, wire336, wire335, wire334, wire333, wire332, wire331, wire330, wire329, wire328, wire327, wire326, wire325, wire324, wire323, wire322, wire321, wire320, wire319, wire318, wire317, wire316, wire315, wire314, wire313, wire312, wire311, wire310, wire309, wire308, wire307, wire306, wire305, wire304, wire303, wire302, wire301, wire300, wire299, wire298, wire297, wire296, wire295, wire294, wire293, wire292, wire291, wire290, wire289, wire288, wire287, wire286, wire285, wire284, wire283, wire282, wire281, wire280, wire279, wire278, wire277, wire276, wire275, wire274, wire273, wire272, wire271, wire270, wire269, wire268, wire267, wire266, wire265, wire264, wire263, wire262, wire261, wire260, wire259, wire258, wire257, wire256, wire255, wire254, wire253, wire252, wire251, wire250, wire249, wire248, wire247, wire246, wire245, wire244, wire243, wire242, wire241, wire240, wire239, wire238, wire237, wire236, wire235, wire234, wire233, wire232, wire231, wire230, wire229, wire228, wire227, wire226, wire225, wire224, wire223, wire222, wire221, wire220, wire219, wire218, wire217, wire216, wire215, wire214, wire213, wire212, wire211, wire210, wire209, wire208, wire207, wire206, wire205, wire204, wire203, wire202, wire201, wire200, wire199, wire198, wire197, wire196, wire195, wire194, wire193, wire192, wire191, wire190, wire189, wire188, wire187, wire186, wire185, wire184, wire183, wire182, wire181, wire180, wire179, wire178, wire177, wire176, wire175, wire174, wire173, wire172, wire171, wire170, wire169, wire168, wire167, wire166, wire165, wire164, wire163, wire162, wire161, wire160, wire159, wire158, wire157, wire156, wire155, wire154, wire153, wire152, wire151, wire150, wire149, wire148, wire147, wire146, wire145, wire144, wire143, wire142, wire141, wire140, wire139, wire138, wire137, wire136, wire135, wire134, wire133, wire132, wire131, wire130, wire129, wire128, wire127, wire126, wire125, wire124, wire123, wire122, wire121, wire120, wire119, wire118, wire117, wire116, wire115, wire114, wire113, wire112, wire111, wire110, wire109, wire108, wire107, wire106, wire105, wire104, wire103, wire102, wire101, wire100, wire99, wire98, wire97, wire96, wire95, wire94, wire93, wire92, wire91, wire90, wire89, wire88, wire87, wire86, wire85, wire84, wire83, wire82, wire81, wire80, wire79, wire78, wire77, wire76, wire75, wire74, wire73, wire72, wire71, wire70, wire69, wire68, wire67, wire66, wire65, wire64, wire63, wire62, wire61, wire60, wire59, wire58, wire57, wire56, wire55, wire54, wire53, wire52, wire51, wire50, wire49, wire48, wire47, wire46, wire45, wire44, wire43, wire42, wire41, wire40, wire39, wire38, wire37, wire36, wire35, wire34, wire33, wire32, wire31, wire30, wire29, wire28, wire27, wire26, wire25, wire24, wire23, wire22, wire21, wire20, wire19, wire18, wire17, wire16, wire15, wire14, wire13, wire12, wire11, wire10, wire9, wire8, wire7, wire6, wire5, wire4, wire3, wire2, wire1, wire0};
    assign out = data_concat;


endmodule

