module select_length(
    input wire [40959:0] data,
    input wire [11:0] sel,
    output wire [9:0] out
);
    wire [4095:0] sel_out;
    select_signal s0(.sel(sel), .out(sel_out));
    muxnm_tristate #(4096, 10) mxt1(.in(data), .sel(sel_out) ,.out(out));

endmodule

module select_signal(
    input wire [11:0] sel,
    output wire [4095:0] out
);
    wire [11:0] buffered_input;
    bufferH4096_12b$ buff(.in(sel), .out(buffered_input));
    equaln #(12) e0(.a(buffered_input), .b(12'b000000000000), .eq(weq0));
    equaln #(12) e1(.a(buffered_input), .b(12'b000000000001), .eq(weq1));
    equaln #(12) e2(.a(buffered_input), .b(12'b000000000010), .eq(weq2));
    equaln #(12) e3(.a(buffered_input), .b(12'b000000000011), .eq(weq3));
    equaln #(12) e4(.a(buffered_input), .b(12'b000000000100), .eq(weq4));
    equaln #(12) e5(.a(buffered_input), .b(12'b000000000101), .eq(weq5));
    equaln #(12) e6(.a(buffered_input), .b(12'b000000000110), .eq(weq6));
    equaln #(12) e7(.a(buffered_input), .b(12'b000000000111), .eq(weq7));
    equaln #(12) e8(.a(buffered_input), .b(12'b000000001000), .eq(weq8));
    equaln #(12) e9(.a(buffered_input), .b(12'b000000001001), .eq(weq9));
    equaln #(12) e10(.a(buffered_input), .b(12'b000000001010), .eq(weq10));
    equaln #(12) e11(.a(buffered_input), .b(12'b000000001011), .eq(weq11));
    equaln #(12) e12(.a(buffered_input), .b(12'b000000001100), .eq(weq12));
    equaln #(12) e13(.a(buffered_input), .b(12'b000000001101), .eq(weq13));
    equaln #(12) e14(.a(buffered_input), .b(12'b000000001110), .eq(weq14));
    equaln #(12) e15(.a(buffered_input), .b(12'b000000001111), .eq(weq15));
    equaln #(12) e16(.a(buffered_input), .b(12'b000000010000), .eq(weq16));
    equaln #(12) e17(.a(buffered_input), .b(12'b000000010001), .eq(weq17));
    equaln #(12) e18(.a(buffered_input), .b(12'b000000010010), .eq(weq18));
    equaln #(12) e19(.a(buffered_input), .b(12'b000000010011), .eq(weq19));
    equaln #(12) e20(.a(buffered_input), .b(12'b000000010100), .eq(weq20));
    equaln #(12) e21(.a(buffered_input), .b(12'b000000010101), .eq(weq21));
    equaln #(12) e22(.a(buffered_input), .b(12'b000000010110), .eq(weq22));
    equaln #(12) e23(.a(buffered_input), .b(12'b000000010111), .eq(weq23));
    equaln #(12) e24(.a(buffered_input), .b(12'b000000011000), .eq(weq24));
    equaln #(12) e25(.a(buffered_input), .b(12'b000000011001), .eq(weq25));
    equaln #(12) e26(.a(buffered_input), .b(12'b000000011010), .eq(weq26));
    equaln #(12) e27(.a(buffered_input), .b(12'b000000011011), .eq(weq27));
    equaln #(12) e28(.a(buffered_input), .b(12'b000000011100), .eq(weq28));
    equaln #(12) e29(.a(buffered_input), .b(12'b000000011101), .eq(weq29));
    equaln #(12) e30(.a(buffered_input), .b(12'b000000011110), .eq(weq30));
    equaln #(12) e31(.a(buffered_input), .b(12'b000000011111), .eq(weq31));
    equaln #(12) e32(.a(buffered_input), .b(12'b000000100000), .eq(weq32));
    equaln #(12) e33(.a(buffered_input), .b(12'b000000100001), .eq(weq33));
    equaln #(12) e34(.a(buffered_input), .b(12'b000000100010), .eq(weq34));
    equaln #(12) e35(.a(buffered_input), .b(12'b000000100011), .eq(weq35));
    equaln #(12) e36(.a(buffered_input), .b(12'b000000100100), .eq(weq36));
    equaln #(12) e37(.a(buffered_input), .b(12'b000000100101), .eq(weq37));
    equaln #(12) e38(.a(buffered_input), .b(12'b000000100110), .eq(weq38));
    equaln #(12) e39(.a(buffered_input), .b(12'b000000100111), .eq(weq39));
    equaln #(12) e40(.a(buffered_input), .b(12'b000000101000), .eq(weq40));
    equaln #(12) e41(.a(buffered_input), .b(12'b000000101001), .eq(weq41));
    equaln #(12) e42(.a(buffered_input), .b(12'b000000101010), .eq(weq42));
    equaln #(12) e43(.a(buffered_input), .b(12'b000000101011), .eq(weq43));
    equaln #(12) e44(.a(buffered_input), .b(12'b000000101100), .eq(weq44));
    equaln #(12) e45(.a(buffered_input), .b(12'b000000101101), .eq(weq45));
    equaln #(12) e46(.a(buffered_input), .b(12'b000000101110), .eq(weq46));
    equaln #(12) e47(.a(buffered_input), .b(12'b000000101111), .eq(weq47));
    equaln #(12) e48(.a(buffered_input), .b(12'b000000110000), .eq(weq48));
    equaln #(12) e49(.a(buffered_input), .b(12'b000000110001), .eq(weq49));
    equaln #(12) e50(.a(buffered_input), .b(12'b000000110010), .eq(weq50));
    equaln #(12) e51(.a(buffered_input), .b(12'b000000110011), .eq(weq51));
    equaln #(12) e52(.a(buffered_input), .b(12'b000000110100), .eq(weq52));
    equaln #(12) e53(.a(buffered_input), .b(12'b000000110101), .eq(weq53));
    equaln #(12) e54(.a(buffered_input), .b(12'b000000110110), .eq(weq54));
    equaln #(12) e55(.a(buffered_input), .b(12'b000000110111), .eq(weq55));
    equaln #(12) e56(.a(buffered_input), .b(12'b000000111000), .eq(weq56));
    equaln #(12) e57(.a(buffered_input), .b(12'b000000111001), .eq(weq57));
    equaln #(12) e58(.a(buffered_input), .b(12'b000000111010), .eq(weq58));
    equaln #(12) e59(.a(buffered_input), .b(12'b000000111011), .eq(weq59));
    equaln #(12) e60(.a(buffered_input), .b(12'b000000111100), .eq(weq60));
    equaln #(12) e61(.a(buffered_input), .b(12'b000000111101), .eq(weq61));
    equaln #(12) e62(.a(buffered_input), .b(12'b000000111110), .eq(weq62));
    equaln #(12) e63(.a(buffered_input), .b(12'b000000111111), .eq(weq63));
    equaln #(12) e64(.a(buffered_input), .b(12'b000001000000), .eq(weq64));
    equaln #(12) e65(.a(buffered_input), .b(12'b000001000001), .eq(weq65));
    equaln #(12) e66(.a(buffered_input), .b(12'b000001000010), .eq(weq66));
    equaln #(12) e67(.a(buffered_input), .b(12'b000001000011), .eq(weq67));
    equaln #(12) e68(.a(buffered_input), .b(12'b000001000100), .eq(weq68));
    equaln #(12) e69(.a(buffered_input), .b(12'b000001000101), .eq(weq69));
    equaln #(12) e70(.a(buffered_input), .b(12'b000001000110), .eq(weq70));
    equaln #(12) e71(.a(buffered_input), .b(12'b000001000111), .eq(weq71));
    equaln #(12) e72(.a(buffered_input), .b(12'b000001001000), .eq(weq72));
    equaln #(12) e73(.a(buffered_input), .b(12'b000001001001), .eq(weq73));
    equaln #(12) e74(.a(buffered_input), .b(12'b000001001010), .eq(weq74));
    equaln #(12) e75(.a(buffered_input), .b(12'b000001001011), .eq(weq75));
    equaln #(12) e76(.a(buffered_input), .b(12'b000001001100), .eq(weq76));
    equaln #(12) e77(.a(buffered_input), .b(12'b000001001101), .eq(weq77));
    equaln #(12) e78(.a(buffered_input), .b(12'b000001001110), .eq(weq78));
    equaln #(12) e79(.a(buffered_input), .b(12'b000001001111), .eq(weq79));
    equaln #(12) e80(.a(buffered_input), .b(12'b000001010000), .eq(weq80));
    equaln #(12) e81(.a(buffered_input), .b(12'b000001010001), .eq(weq81));
    equaln #(12) e82(.a(buffered_input), .b(12'b000001010010), .eq(weq82));
    equaln #(12) e83(.a(buffered_input), .b(12'b000001010011), .eq(weq83));
    equaln #(12) e84(.a(buffered_input), .b(12'b000001010100), .eq(weq84));
    equaln #(12) e85(.a(buffered_input), .b(12'b000001010101), .eq(weq85));
    equaln #(12) e86(.a(buffered_input), .b(12'b000001010110), .eq(weq86));
    equaln #(12) e87(.a(buffered_input), .b(12'b000001010111), .eq(weq87));
    equaln #(12) e88(.a(buffered_input), .b(12'b000001011000), .eq(weq88));
    equaln #(12) e89(.a(buffered_input), .b(12'b000001011001), .eq(weq89));
    equaln #(12) e90(.a(buffered_input), .b(12'b000001011010), .eq(weq90));
    equaln #(12) e91(.a(buffered_input), .b(12'b000001011011), .eq(weq91));
    equaln #(12) e92(.a(buffered_input), .b(12'b000001011100), .eq(weq92));
    equaln #(12) e93(.a(buffered_input), .b(12'b000001011101), .eq(weq93));
    equaln #(12) e94(.a(buffered_input), .b(12'b000001011110), .eq(weq94));
    equaln #(12) e95(.a(buffered_input), .b(12'b000001011111), .eq(weq95));
    equaln #(12) e96(.a(buffered_input), .b(12'b000001100000), .eq(weq96));
    equaln #(12) e97(.a(buffered_input), .b(12'b000001100001), .eq(weq97));
    equaln #(12) e98(.a(buffered_input), .b(12'b000001100010), .eq(weq98));
    equaln #(12) e99(.a(buffered_input), .b(12'b000001100011), .eq(weq99));
    equaln #(12) e100(.a(buffered_input), .b(12'b000001100100), .eq(weq100));
    equaln #(12) e101(.a(buffered_input), .b(12'b000001100101), .eq(weq101));
    equaln #(12) e102(.a(buffered_input), .b(12'b000001100110), .eq(weq102));
    equaln #(12) e103(.a(buffered_input), .b(12'b000001100111), .eq(weq103));
    equaln #(12) e104(.a(buffered_input), .b(12'b000001101000), .eq(weq104));
    equaln #(12) e105(.a(buffered_input), .b(12'b000001101001), .eq(weq105));
    equaln #(12) e106(.a(buffered_input), .b(12'b000001101010), .eq(weq106));
    equaln #(12) e107(.a(buffered_input), .b(12'b000001101011), .eq(weq107));
    equaln #(12) e108(.a(buffered_input), .b(12'b000001101100), .eq(weq108));
    equaln #(12) e109(.a(buffered_input), .b(12'b000001101101), .eq(weq109));
    equaln #(12) e110(.a(buffered_input), .b(12'b000001101110), .eq(weq110));
    equaln #(12) e111(.a(buffered_input), .b(12'b000001101111), .eq(weq111));
    equaln #(12) e112(.a(buffered_input), .b(12'b000001110000), .eq(weq112));
    equaln #(12) e113(.a(buffered_input), .b(12'b000001110001), .eq(weq113));
    equaln #(12) e114(.a(buffered_input), .b(12'b000001110010), .eq(weq114));
    equaln #(12) e115(.a(buffered_input), .b(12'b000001110011), .eq(weq115));
    equaln #(12) e116(.a(buffered_input), .b(12'b000001110100), .eq(weq116));
    equaln #(12) e117(.a(buffered_input), .b(12'b000001110101), .eq(weq117));
    equaln #(12) e118(.a(buffered_input), .b(12'b000001110110), .eq(weq118));
    equaln #(12) e119(.a(buffered_input), .b(12'b000001110111), .eq(weq119));
    equaln #(12) e120(.a(buffered_input), .b(12'b000001111000), .eq(weq120));
    equaln #(12) e121(.a(buffered_input), .b(12'b000001111001), .eq(weq121));
    equaln #(12) e122(.a(buffered_input), .b(12'b000001111010), .eq(weq122));
    equaln #(12) e123(.a(buffered_input), .b(12'b000001111011), .eq(weq123));
    equaln #(12) e124(.a(buffered_input), .b(12'b000001111100), .eq(weq124));
    equaln #(12) e125(.a(buffered_input), .b(12'b000001111101), .eq(weq125));
    equaln #(12) e126(.a(buffered_input), .b(12'b000001111110), .eq(weq126));
    equaln #(12) e127(.a(buffered_input), .b(12'b000001111111), .eq(weq127));
    equaln #(12) e128(.a(buffered_input), .b(12'b000010000000), .eq(weq128));
    equaln #(12) e129(.a(buffered_input), .b(12'b000010000001), .eq(weq129));
    equaln #(12) e130(.a(buffered_input), .b(12'b000010000010), .eq(weq130));
    equaln #(12) e131(.a(buffered_input), .b(12'b000010000011), .eq(weq131));
    equaln #(12) e132(.a(buffered_input), .b(12'b000010000100), .eq(weq132));
    equaln #(12) e133(.a(buffered_input), .b(12'b000010000101), .eq(weq133));
    equaln #(12) e134(.a(buffered_input), .b(12'b000010000110), .eq(weq134));
    equaln #(12) e135(.a(buffered_input), .b(12'b000010000111), .eq(weq135));
    equaln #(12) e136(.a(buffered_input), .b(12'b000010001000), .eq(weq136));
    equaln #(12) e137(.a(buffered_input), .b(12'b000010001001), .eq(weq137));
    equaln #(12) e138(.a(buffered_input), .b(12'b000010001010), .eq(weq138));
    equaln #(12) e139(.a(buffered_input), .b(12'b000010001011), .eq(weq139));
    equaln #(12) e140(.a(buffered_input), .b(12'b000010001100), .eq(weq140));
    equaln #(12) e141(.a(buffered_input), .b(12'b000010001101), .eq(weq141));
    equaln #(12) e142(.a(buffered_input), .b(12'b000010001110), .eq(weq142));
    equaln #(12) e143(.a(buffered_input), .b(12'b000010001111), .eq(weq143));
    equaln #(12) e144(.a(buffered_input), .b(12'b000010010000), .eq(weq144));
    equaln #(12) e145(.a(buffered_input), .b(12'b000010010001), .eq(weq145));
    equaln #(12) e146(.a(buffered_input), .b(12'b000010010010), .eq(weq146));
    equaln #(12) e147(.a(buffered_input), .b(12'b000010010011), .eq(weq147));
    equaln #(12) e148(.a(buffered_input), .b(12'b000010010100), .eq(weq148));
    equaln #(12) e149(.a(buffered_input), .b(12'b000010010101), .eq(weq149));
    equaln #(12) e150(.a(buffered_input), .b(12'b000010010110), .eq(weq150));
    equaln #(12) e151(.a(buffered_input), .b(12'b000010010111), .eq(weq151));
    equaln #(12) e152(.a(buffered_input), .b(12'b000010011000), .eq(weq152));
    equaln #(12) e153(.a(buffered_input), .b(12'b000010011001), .eq(weq153));
    equaln #(12) e154(.a(buffered_input), .b(12'b000010011010), .eq(weq154));
    equaln #(12) e155(.a(buffered_input), .b(12'b000010011011), .eq(weq155));
    equaln #(12) e156(.a(buffered_input), .b(12'b000010011100), .eq(weq156));
    equaln #(12) e157(.a(buffered_input), .b(12'b000010011101), .eq(weq157));
    equaln #(12) e158(.a(buffered_input), .b(12'b000010011110), .eq(weq158));
    equaln #(12) e159(.a(buffered_input), .b(12'b000010011111), .eq(weq159));
    equaln #(12) e160(.a(buffered_input), .b(12'b000010100000), .eq(weq160));
    equaln #(12) e161(.a(buffered_input), .b(12'b000010100001), .eq(weq161));
    equaln #(12) e162(.a(buffered_input), .b(12'b000010100010), .eq(weq162));
    equaln #(12) e163(.a(buffered_input), .b(12'b000010100011), .eq(weq163));
    equaln #(12) e164(.a(buffered_input), .b(12'b000010100100), .eq(weq164));
    equaln #(12) e165(.a(buffered_input), .b(12'b000010100101), .eq(weq165));
    equaln #(12) e166(.a(buffered_input), .b(12'b000010100110), .eq(weq166));
    equaln #(12) e167(.a(buffered_input), .b(12'b000010100111), .eq(weq167));
    equaln #(12) e168(.a(buffered_input), .b(12'b000010101000), .eq(weq168));
    equaln #(12) e169(.a(buffered_input), .b(12'b000010101001), .eq(weq169));
    equaln #(12) e170(.a(buffered_input), .b(12'b000010101010), .eq(weq170));
    equaln #(12) e171(.a(buffered_input), .b(12'b000010101011), .eq(weq171));
    equaln #(12) e172(.a(buffered_input), .b(12'b000010101100), .eq(weq172));
    equaln #(12) e173(.a(buffered_input), .b(12'b000010101101), .eq(weq173));
    equaln #(12) e174(.a(buffered_input), .b(12'b000010101110), .eq(weq174));
    equaln #(12) e175(.a(buffered_input), .b(12'b000010101111), .eq(weq175));
    equaln #(12) e176(.a(buffered_input), .b(12'b000010110000), .eq(weq176));
    equaln #(12) e177(.a(buffered_input), .b(12'b000010110001), .eq(weq177));
    equaln #(12) e178(.a(buffered_input), .b(12'b000010110010), .eq(weq178));
    equaln #(12) e179(.a(buffered_input), .b(12'b000010110011), .eq(weq179));
    equaln #(12) e180(.a(buffered_input), .b(12'b000010110100), .eq(weq180));
    equaln #(12) e181(.a(buffered_input), .b(12'b000010110101), .eq(weq181));
    equaln #(12) e182(.a(buffered_input), .b(12'b000010110110), .eq(weq182));
    equaln #(12) e183(.a(buffered_input), .b(12'b000010110111), .eq(weq183));
    equaln #(12) e184(.a(buffered_input), .b(12'b000010111000), .eq(weq184));
    equaln #(12) e185(.a(buffered_input), .b(12'b000010111001), .eq(weq185));
    equaln #(12) e186(.a(buffered_input), .b(12'b000010111010), .eq(weq186));
    equaln #(12) e187(.a(buffered_input), .b(12'b000010111011), .eq(weq187));
    equaln #(12) e188(.a(buffered_input), .b(12'b000010111100), .eq(weq188));
    equaln #(12) e189(.a(buffered_input), .b(12'b000010111101), .eq(weq189));
    equaln #(12) e190(.a(buffered_input), .b(12'b000010111110), .eq(weq190));
    equaln #(12) e191(.a(buffered_input), .b(12'b000010111111), .eq(weq191));
    equaln #(12) e192(.a(buffered_input), .b(12'b000011000000), .eq(weq192));
    equaln #(12) e193(.a(buffered_input), .b(12'b000011000001), .eq(weq193));
    equaln #(12) e194(.a(buffered_input), .b(12'b000011000010), .eq(weq194));
    equaln #(12) e195(.a(buffered_input), .b(12'b000011000011), .eq(weq195));
    equaln #(12) e196(.a(buffered_input), .b(12'b000011000100), .eq(weq196));
    equaln #(12) e197(.a(buffered_input), .b(12'b000011000101), .eq(weq197));
    equaln #(12) e198(.a(buffered_input), .b(12'b000011000110), .eq(weq198));
    equaln #(12) e199(.a(buffered_input), .b(12'b000011000111), .eq(weq199));
    equaln #(12) e200(.a(buffered_input), .b(12'b000011001000), .eq(weq200));
    equaln #(12) e201(.a(buffered_input), .b(12'b000011001001), .eq(weq201));
    equaln #(12) e202(.a(buffered_input), .b(12'b000011001010), .eq(weq202));
    equaln #(12) e203(.a(buffered_input), .b(12'b000011001011), .eq(weq203));
    equaln #(12) e204(.a(buffered_input), .b(12'b000011001100), .eq(weq204));
    equaln #(12) e205(.a(buffered_input), .b(12'b000011001101), .eq(weq205));
    equaln #(12) e206(.a(buffered_input), .b(12'b000011001110), .eq(weq206));
    equaln #(12) e207(.a(buffered_input), .b(12'b000011001111), .eq(weq207));
    equaln #(12) e208(.a(buffered_input), .b(12'b000011010000), .eq(weq208));
    equaln #(12) e209(.a(buffered_input), .b(12'b000011010001), .eq(weq209));
    equaln #(12) e210(.a(buffered_input), .b(12'b000011010010), .eq(weq210));
    equaln #(12) e211(.a(buffered_input), .b(12'b000011010011), .eq(weq211));
    equaln #(12) e212(.a(buffered_input), .b(12'b000011010100), .eq(weq212));
    equaln #(12) e213(.a(buffered_input), .b(12'b000011010101), .eq(weq213));
    equaln #(12) e214(.a(buffered_input), .b(12'b000011010110), .eq(weq214));
    equaln #(12) e215(.a(buffered_input), .b(12'b000011010111), .eq(weq215));
    equaln #(12) e216(.a(buffered_input), .b(12'b000011011000), .eq(weq216));
    equaln #(12) e217(.a(buffered_input), .b(12'b000011011001), .eq(weq217));
    equaln #(12) e218(.a(buffered_input), .b(12'b000011011010), .eq(weq218));
    equaln #(12) e219(.a(buffered_input), .b(12'b000011011011), .eq(weq219));
    equaln #(12) e220(.a(buffered_input), .b(12'b000011011100), .eq(weq220));
    equaln #(12) e221(.a(buffered_input), .b(12'b000011011101), .eq(weq221));
    equaln #(12) e222(.a(buffered_input), .b(12'b000011011110), .eq(weq222));
    equaln #(12) e223(.a(buffered_input), .b(12'b000011011111), .eq(weq223));
    equaln #(12) e224(.a(buffered_input), .b(12'b000011100000), .eq(weq224));
    equaln #(12) e225(.a(buffered_input), .b(12'b000011100001), .eq(weq225));
    equaln #(12) e226(.a(buffered_input), .b(12'b000011100010), .eq(weq226));
    equaln #(12) e227(.a(buffered_input), .b(12'b000011100011), .eq(weq227));
    equaln #(12) e228(.a(buffered_input), .b(12'b000011100100), .eq(weq228));
    equaln #(12) e229(.a(buffered_input), .b(12'b000011100101), .eq(weq229));
    equaln #(12) e230(.a(buffered_input), .b(12'b000011100110), .eq(weq230));
    equaln #(12) e231(.a(buffered_input), .b(12'b000011100111), .eq(weq231));
    equaln #(12) e232(.a(buffered_input), .b(12'b000011101000), .eq(weq232));
    equaln #(12) e233(.a(buffered_input), .b(12'b000011101001), .eq(weq233));
    equaln #(12) e234(.a(buffered_input), .b(12'b000011101010), .eq(weq234));
    equaln #(12) e235(.a(buffered_input), .b(12'b000011101011), .eq(weq235));
    equaln #(12) e236(.a(buffered_input), .b(12'b000011101100), .eq(weq236));
    equaln #(12) e237(.a(buffered_input), .b(12'b000011101101), .eq(weq237));
    equaln #(12) e238(.a(buffered_input), .b(12'b000011101110), .eq(weq238));
    equaln #(12) e239(.a(buffered_input), .b(12'b000011101111), .eq(weq239));
    equaln #(12) e240(.a(buffered_input), .b(12'b000011110000), .eq(weq240));
    equaln #(12) e241(.a(buffered_input), .b(12'b000011110001), .eq(weq241));
    equaln #(12) e242(.a(buffered_input), .b(12'b000011110010), .eq(weq242));
    equaln #(12) e243(.a(buffered_input), .b(12'b000011110011), .eq(weq243));
    equaln #(12) e244(.a(buffered_input), .b(12'b000011110100), .eq(weq244));
    equaln #(12) e245(.a(buffered_input), .b(12'b000011110101), .eq(weq245));
    equaln #(12) e246(.a(buffered_input), .b(12'b000011110110), .eq(weq246));
    equaln #(12) e247(.a(buffered_input), .b(12'b000011110111), .eq(weq247));
    equaln #(12) e248(.a(buffered_input), .b(12'b000011111000), .eq(weq248));
    equaln #(12) e249(.a(buffered_input), .b(12'b000011111001), .eq(weq249));
    equaln #(12) e250(.a(buffered_input), .b(12'b000011111010), .eq(weq250));
    equaln #(12) e251(.a(buffered_input), .b(12'b000011111011), .eq(weq251));
    equaln #(12) e252(.a(buffered_input), .b(12'b000011111100), .eq(weq252));
    equaln #(12) e253(.a(buffered_input), .b(12'b000011111101), .eq(weq253));
    equaln #(12) e254(.a(buffered_input), .b(12'b000011111110), .eq(weq254));
    equaln #(12) e255(.a(buffered_input), .b(12'b000011111111), .eq(weq255));
    equaln #(12) e256(.a(buffered_input), .b(12'b000100000000), .eq(weq256));
    equaln #(12) e257(.a(buffered_input), .b(12'b000100000001), .eq(weq257));
    equaln #(12) e258(.a(buffered_input), .b(12'b000100000010), .eq(weq258));
    equaln #(12) e259(.a(buffered_input), .b(12'b000100000011), .eq(weq259));
    equaln #(12) e260(.a(buffered_input), .b(12'b000100000100), .eq(weq260));
    equaln #(12) e261(.a(buffered_input), .b(12'b000100000101), .eq(weq261));
    equaln #(12) e262(.a(buffered_input), .b(12'b000100000110), .eq(weq262));
    equaln #(12) e263(.a(buffered_input), .b(12'b000100000111), .eq(weq263));
    equaln #(12) e264(.a(buffered_input), .b(12'b000100001000), .eq(weq264));
    equaln #(12) e265(.a(buffered_input), .b(12'b000100001001), .eq(weq265));
    equaln #(12) e266(.a(buffered_input), .b(12'b000100001010), .eq(weq266));
    equaln #(12) e267(.a(buffered_input), .b(12'b000100001011), .eq(weq267));
    equaln #(12) e268(.a(buffered_input), .b(12'b000100001100), .eq(weq268));
    equaln #(12) e269(.a(buffered_input), .b(12'b000100001101), .eq(weq269));
    equaln #(12) e270(.a(buffered_input), .b(12'b000100001110), .eq(weq270));
    equaln #(12) e271(.a(buffered_input), .b(12'b000100001111), .eq(weq271));
    equaln #(12) e272(.a(buffered_input), .b(12'b000100010000), .eq(weq272));
    equaln #(12) e273(.a(buffered_input), .b(12'b000100010001), .eq(weq273));
    equaln #(12) e274(.a(buffered_input), .b(12'b000100010010), .eq(weq274));
    equaln #(12) e275(.a(buffered_input), .b(12'b000100010011), .eq(weq275));
    equaln #(12) e276(.a(buffered_input), .b(12'b000100010100), .eq(weq276));
    equaln #(12) e277(.a(buffered_input), .b(12'b000100010101), .eq(weq277));
    equaln #(12) e278(.a(buffered_input), .b(12'b000100010110), .eq(weq278));
    equaln #(12) e279(.a(buffered_input), .b(12'b000100010111), .eq(weq279));
    equaln #(12) e280(.a(buffered_input), .b(12'b000100011000), .eq(weq280));
    equaln #(12) e281(.a(buffered_input), .b(12'b000100011001), .eq(weq281));
    equaln #(12) e282(.a(buffered_input), .b(12'b000100011010), .eq(weq282));
    equaln #(12) e283(.a(buffered_input), .b(12'b000100011011), .eq(weq283));
    equaln #(12) e284(.a(buffered_input), .b(12'b000100011100), .eq(weq284));
    equaln #(12) e285(.a(buffered_input), .b(12'b000100011101), .eq(weq285));
    equaln #(12) e286(.a(buffered_input), .b(12'b000100011110), .eq(weq286));
    equaln #(12) e287(.a(buffered_input), .b(12'b000100011111), .eq(weq287));
    equaln #(12) e288(.a(buffered_input), .b(12'b000100100000), .eq(weq288));
    equaln #(12) e289(.a(buffered_input), .b(12'b000100100001), .eq(weq289));
    equaln #(12) e290(.a(buffered_input), .b(12'b000100100010), .eq(weq290));
    equaln #(12) e291(.a(buffered_input), .b(12'b000100100011), .eq(weq291));
    equaln #(12) e292(.a(buffered_input), .b(12'b000100100100), .eq(weq292));
    equaln #(12) e293(.a(buffered_input), .b(12'b000100100101), .eq(weq293));
    equaln #(12) e294(.a(buffered_input), .b(12'b000100100110), .eq(weq294));
    equaln #(12) e295(.a(buffered_input), .b(12'b000100100111), .eq(weq295));
    equaln #(12) e296(.a(buffered_input), .b(12'b000100101000), .eq(weq296));
    equaln #(12) e297(.a(buffered_input), .b(12'b000100101001), .eq(weq297));
    equaln #(12) e298(.a(buffered_input), .b(12'b000100101010), .eq(weq298));
    equaln #(12) e299(.a(buffered_input), .b(12'b000100101011), .eq(weq299));
    equaln #(12) e300(.a(buffered_input), .b(12'b000100101100), .eq(weq300));
    equaln #(12) e301(.a(buffered_input), .b(12'b000100101101), .eq(weq301));
    equaln #(12) e302(.a(buffered_input), .b(12'b000100101110), .eq(weq302));
    equaln #(12) e303(.a(buffered_input), .b(12'b000100101111), .eq(weq303));
    equaln #(12) e304(.a(buffered_input), .b(12'b000100110000), .eq(weq304));
    equaln #(12) e305(.a(buffered_input), .b(12'b000100110001), .eq(weq305));
    equaln #(12) e306(.a(buffered_input), .b(12'b000100110010), .eq(weq306));
    equaln #(12) e307(.a(buffered_input), .b(12'b000100110011), .eq(weq307));
    equaln #(12) e308(.a(buffered_input), .b(12'b000100110100), .eq(weq308));
    equaln #(12) e309(.a(buffered_input), .b(12'b000100110101), .eq(weq309));
    equaln #(12) e310(.a(buffered_input), .b(12'b000100110110), .eq(weq310));
    equaln #(12) e311(.a(buffered_input), .b(12'b000100110111), .eq(weq311));
    equaln #(12) e312(.a(buffered_input), .b(12'b000100111000), .eq(weq312));
    equaln #(12) e313(.a(buffered_input), .b(12'b000100111001), .eq(weq313));
    equaln #(12) e314(.a(buffered_input), .b(12'b000100111010), .eq(weq314));
    equaln #(12) e315(.a(buffered_input), .b(12'b000100111011), .eq(weq315));
    equaln #(12) e316(.a(buffered_input), .b(12'b000100111100), .eq(weq316));
    equaln #(12) e317(.a(buffered_input), .b(12'b000100111101), .eq(weq317));
    equaln #(12) e318(.a(buffered_input), .b(12'b000100111110), .eq(weq318));
    equaln #(12) e319(.a(buffered_input), .b(12'b000100111111), .eq(weq319));
    equaln #(12) e320(.a(buffered_input), .b(12'b000101000000), .eq(weq320));
    equaln #(12) e321(.a(buffered_input), .b(12'b000101000001), .eq(weq321));
    equaln #(12) e322(.a(buffered_input), .b(12'b000101000010), .eq(weq322));
    equaln #(12) e323(.a(buffered_input), .b(12'b000101000011), .eq(weq323));
    equaln #(12) e324(.a(buffered_input), .b(12'b000101000100), .eq(weq324));
    equaln #(12) e325(.a(buffered_input), .b(12'b000101000101), .eq(weq325));
    equaln #(12) e326(.a(buffered_input), .b(12'b000101000110), .eq(weq326));
    equaln #(12) e327(.a(buffered_input), .b(12'b000101000111), .eq(weq327));
    equaln #(12) e328(.a(buffered_input), .b(12'b000101001000), .eq(weq328));
    equaln #(12) e329(.a(buffered_input), .b(12'b000101001001), .eq(weq329));
    equaln #(12) e330(.a(buffered_input), .b(12'b000101001010), .eq(weq330));
    equaln #(12) e331(.a(buffered_input), .b(12'b000101001011), .eq(weq331));
    equaln #(12) e332(.a(buffered_input), .b(12'b000101001100), .eq(weq332));
    equaln #(12) e333(.a(buffered_input), .b(12'b000101001101), .eq(weq333));
    equaln #(12) e334(.a(buffered_input), .b(12'b000101001110), .eq(weq334));
    equaln #(12) e335(.a(buffered_input), .b(12'b000101001111), .eq(weq335));
    equaln #(12) e336(.a(buffered_input), .b(12'b000101010000), .eq(weq336));
    equaln #(12) e337(.a(buffered_input), .b(12'b000101010001), .eq(weq337));
    equaln #(12) e338(.a(buffered_input), .b(12'b000101010010), .eq(weq338));
    equaln #(12) e339(.a(buffered_input), .b(12'b000101010011), .eq(weq339));
    equaln #(12) e340(.a(buffered_input), .b(12'b000101010100), .eq(weq340));
    equaln #(12) e341(.a(buffered_input), .b(12'b000101010101), .eq(weq341));
    equaln #(12) e342(.a(buffered_input), .b(12'b000101010110), .eq(weq342));
    equaln #(12) e343(.a(buffered_input), .b(12'b000101010111), .eq(weq343));
    equaln #(12) e344(.a(buffered_input), .b(12'b000101011000), .eq(weq344));
    equaln #(12) e345(.a(buffered_input), .b(12'b000101011001), .eq(weq345));
    equaln #(12) e346(.a(buffered_input), .b(12'b000101011010), .eq(weq346));
    equaln #(12) e347(.a(buffered_input), .b(12'b000101011011), .eq(weq347));
    equaln #(12) e348(.a(buffered_input), .b(12'b000101011100), .eq(weq348));
    equaln #(12) e349(.a(buffered_input), .b(12'b000101011101), .eq(weq349));
    equaln #(12) e350(.a(buffered_input), .b(12'b000101011110), .eq(weq350));
    equaln #(12) e351(.a(buffered_input), .b(12'b000101011111), .eq(weq351));
    equaln #(12) e352(.a(buffered_input), .b(12'b000101100000), .eq(weq352));
    equaln #(12) e353(.a(buffered_input), .b(12'b000101100001), .eq(weq353));
    equaln #(12) e354(.a(buffered_input), .b(12'b000101100010), .eq(weq354));
    equaln #(12) e355(.a(buffered_input), .b(12'b000101100011), .eq(weq355));
    equaln #(12) e356(.a(buffered_input), .b(12'b000101100100), .eq(weq356));
    equaln #(12) e357(.a(buffered_input), .b(12'b000101100101), .eq(weq357));
    equaln #(12) e358(.a(buffered_input), .b(12'b000101100110), .eq(weq358));
    equaln #(12) e359(.a(buffered_input), .b(12'b000101100111), .eq(weq359));
    equaln #(12) e360(.a(buffered_input), .b(12'b000101101000), .eq(weq360));
    equaln #(12) e361(.a(buffered_input), .b(12'b000101101001), .eq(weq361));
    equaln #(12) e362(.a(buffered_input), .b(12'b000101101010), .eq(weq362));
    equaln #(12) e363(.a(buffered_input), .b(12'b000101101011), .eq(weq363));
    equaln #(12) e364(.a(buffered_input), .b(12'b000101101100), .eq(weq364));
    equaln #(12) e365(.a(buffered_input), .b(12'b000101101101), .eq(weq365));
    equaln #(12) e366(.a(buffered_input), .b(12'b000101101110), .eq(weq366));
    equaln #(12) e367(.a(buffered_input), .b(12'b000101101111), .eq(weq367));
    equaln #(12) e368(.a(buffered_input), .b(12'b000101110000), .eq(weq368));
    equaln #(12) e369(.a(buffered_input), .b(12'b000101110001), .eq(weq369));
    equaln #(12) e370(.a(buffered_input), .b(12'b000101110010), .eq(weq370));
    equaln #(12) e371(.a(buffered_input), .b(12'b000101110011), .eq(weq371));
    equaln #(12) e372(.a(buffered_input), .b(12'b000101110100), .eq(weq372));
    equaln #(12) e373(.a(buffered_input), .b(12'b000101110101), .eq(weq373));
    equaln #(12) e374(.a(buffered_input), .b(12'b000101110110), .eq(weq374));
    equaln #(12) e375(.a(buffered_input), .b(12'b000101110111), .eq(weq375));
    equaln #(12) e376(.a(buffered_input), .b(12'b000101111000), .eq(weq376));
    equaln #(12) e377(.a(buffered_input), .b(12'b000101111001), .eq(weq377));
    equaln #(12) e378(.a(buffered_input), .b(12'b000101111010), .eq(weq378));
    equaln #(12) e379(.a(buffered_input), .b(12'b000101111011), .eq(weq379));
    equaln #(12) e380(.a(buffered_input), .b(12'b000101111100), .eq(weq380));
    equaln #(12) e381(.a(buffered_input), .b(12'b000101111101), .eq(weq381));
    equaln #(12) e382(.a(buffered_input), .b(12'b000101111110), .eq(weq382));
    equaln #(12) e383(.a(buffered_input), .b(12'b000101111111), .eq(weq383));
    equaln #(12) e384(.a(buffered_input), .b(12'b000110000000), .eq(weq384));
    equaln #(12) e385(.a(buffered_input), .b(12'b000110000001), .eq(weq385));
    equaln #(12) e386(.a(buffered_input), .b(12'b000110000010), .eq(weq386));
    equaln #(12) e387(.a(buffered_input), .b(12'b000110000011), .eq(weq387));
    equaln #(12) e388(.a(buffered_input), .b(12'b000110000100), .eq(weq388));
    equaln #(12) e389(.a(buffered_input), .b(12'b000110000101), .eq(weq389));
    equaln #(12) e390(.a(buffered_input), .b(12'b000110000110), .eq(weq390));
    equaln #(12) e391(.a(buffered_input), .b(12'b000110000111), .eq(weq391));
    equaln #(12) e392(.a(buffered_input), .b(12'b000110001000), .eq(weq392));
    equaln #(12) e393(.a(buffered_input), .b(12'b000110001001), .eq(weq393));
    equaln #(12) e394(.a(buffered_input), .b(12'b000110001010), .eq(weq394));
    equaln #(12) e395(.a(buffered_input), .b(12'b000110001011), .eq(weq395));
    equaln #(12) e396(.a(buffered_input), .b(12'b000110001100), .eq(weq396));
    equaln #(12) e397(.a(buffered_input), .b(12'b000110001101), .eq(weq397));
    equaln #(12) e398(.a(buffered_input), .b(12'b000110001110), .eq(weq398));
    equaln #(12) e399(.a(buffered_input), .b(12'b000110001111), .eq(weq399));
    equaln #(12) e400(.a(buffered_input), .b(12'b000110010000), .eq(weq400));
    equaln #(12) e401(.a(buffered_input), .b(12'b000110010001), .eq(weq401));
    equaln #(12) e402(.a(buffered_input), .b(12'b000110010010), .eq(weq402));
    equaln #(12) e403(.a(buffered_input), .b(12'b000110010011), .eq(weq403));
    equaln #(12) e404(.a(buffered_input), .b(12'b000110010100), .eq(weq404));
    equaln #(12) e405(.a(buffered_input), .b(12'b000110010101), .eq(weq405));
    equaln #(12) e406(.a(buffered_input), .b(12'b000110010110), .eq(weq406));
    equaln #(12) e407(.a(buffered_input), .b(12'b000110010111), .eq(weq407));
    equaln #(12) e408(.a(buffered_input), .b(12'b000110011000), .eq(weq408));
    equaln #(12) e409(.a(buffered_input), .b(12'b000110011001), .eq(weq409));
    equaln #(12) e410(.a(buffered_input), .b(12'b000110011010), .eq(weq410));
    equaln #(12) e411(.a(buffered_input), .b(12'b000110011011), .eq(weq411));
    equaln #(12) e412(.a(buffered_input), .b(12'b000110011100), .eq(weq412));
    equaln #(12) e413(.a(buffered_input), .b(12'b000110011101), .eq(weq413));
    equaln #(12) e414(.a(buffered_input), .b(12'b000110011110), .eq(weq414));
    equaln #(12) e415(.a(buffered_input), .b(12'b000110011111), .eq(weq415));
    equaln #(12) e416(.a(buffered_input), .b(12'b000110100000), .eq(weq416));
    equaln #(12) e417(.a(buffered_input), .b(12'b000110100001), .eq(weq417));
    equaln #(12) e418(.a(buffered_input), .b(12'b000110100010), .eq(weq418));
    equaln #(12) e419(.a(buffered_input), .b(12'b000110100011), .eq(weq419));
    equaln #(12) e420(.a(buffered_input), .b(12'b000110100100), .eq(weq420));
    equaln #(12) e421(.a(buffered_input), .b(12'b000110100101), .eq(weq421));
    equaln #(12) e422(.a(buffered_input), .b(12'b000110100110), .eq(weq422));
    equaln #(12) e423(.a(buffered_input), .b(12'b000110100111), .eq(weq423));
    equaln #(12) e424(.a(buffered_input), .b(12'b000110101000), .eq(weq424));
    equaln #(12) e425(.a(buffered_input), .b(12'b000110101001), .eq(weq425));
    equaln #(12) e426(.a(buffered_input), .b(12'b000110101010), .eq(weq426));
    equaln #(12) e427(.a(buffered_input), .b(12'b000110101011), .eq(weq427));
    equaln #(12) e428(.a(buffered_input), .b(12'b000110101100), .eq(weq428));
    equaln #(12) e429(.a(buffered_input), .b(12'b000110101101), .eq(weq429));
    equaln #(12) e430(.a(buffered_input), .b(12'b000110101110), .eq(weq430));
    equaln #(12) e431(.a(buffered_input), .b(12'b000110101111), .eq(weq431));
    equaln #(12) e432(.a(buffered_input), .b(12'b000110110000), .eq(weq432));
    equaln #(12) e433(.a(buffered_input), .b(12'b000110110001), .eq(weq433));
    equaln #(12) e434(.a(buffered_input), .b(12'b000110110010), .eq(weq434));
    equaln #(12) e435(.a(buffered_input), .b(12'b000110110011), .eq(weq435));
    equaln #(12) e436(.a(buffered_input), .b(12'b000110110100), .eq(weq436));
    equaln #(12) e437(.a(buffered_input), .b(12'b000110110101), .eq(weq437));
    equaln #(12) e438(.a(buffered_input), .b(12'b000110110110), .eq(weq438));
    equaln #(12) e439(.a(buffered_input), .b(12'b000110110111), .eq(weq439));
    equaln #(12) e440(.a(buffered_input), .b(12'b000110111000), .eq(weq440));
    equaln #(12) e441(.a(buffered_input), .b(12'b000110111001), .eq(weq441));
    equaln #(12) e442(.a(buffered_input), .b(12'b000110111010), .eq(weq442));
    equaln #(12) e443(.a(buffered_input), .b(12'b000110111011), .eq(weq443));
    equaln #(12) e444(.a(buffered_input), .b(12'b000110111100), .eq(weq444));
    equaln #(12) e445(.a(buffered_input), .b(12'b000110111101), .eq(weq445));
    equaln #(12) e446(.a(buffered_input), .b(12'b000110111110), .eq(weq446));
    equaln #(12) e447(.a(buffered_input), .b(12'b000110111111), .eq(weq447));
    equaln #(12) e448(.a(buffered_input), .b(12'b000111000000), .eq(weq448));
    equaln #(12) e449(.a(buffered_input), .b(12'b000111000001), .eq(weq449));
    equaln #(12) e450(.a(buffered_input), .b(12'b000111000010), .eq(weq450));
    equaln #(12) e451(.a(buffered_input), .b(12'b000111000011), .eq(weq451));
    equaln #(12) e452(.a(buffered_input), .b(12'b000111000100), .eq(weq452));
    equaln #(12) e453(.a(buffered_input), .b(12'b000111000101), .eq(weq453));
    equaln #(12) e454(.a(buffered_input), .b(12'b000111000110), .eq(weq454));
    equaln #(12) e455(.a(buffered_input), .b(12'b000111000111), .eq(weq455));
    equaln #(12) e456(.a(buffered_input), .b(12'b000111001000), .eq(weq456));
    equaln #(12) e457(.a(buffered_input), .b(12'b000111001001), .eq(weq457));
    equaln #(12) e458(.a(buffered_input), .b(12'b000111001010), .eq(weq458));
    equaln #(12) e459(.a(buffered_input), .b(12'b000111001011), .eq(weq459));
    equaln #(12) e460(.a(buffered_input), .b(12'b000111001100), .eq(weq460));
    equaln #(12) e461(.a(buffered_input), .b(12'b000111001101), .eq(weq461));
    equaln #(12) e462(.a(buffered_input), .b(12'b000111001110), .eq(weq462));
    equaln #(12) e463(.a(buffered_input), .b(12'b000111001111), .eq(weq463));
    equaln #(12) e464(.a(buffered_input), .b(12'b000111010000), .eq(weq464));
    equaln #(12) e465(.a(buffered_input), .b(12'b000111010001), .eq(weq465));
    equaln #(12) e466(.a(buffered_input), .b(12'b000111010010), .eq(weq466));
    equaln #(12) e467(.a(buffered_input), .b(12'b000111010011), .eq(weq467));
    equaln #(12) e468(.a(buffered_input), .b(12'b000111010100), .eq(weq468));
    equaln #(12) e469(.a(buffered_input), .b(12'b000111010101), .eq(weq469));
    equaln #(12) e470(.a(buffered_input), .b(12'b000111010110), .eq(weq470));
    equaln #(12) e471(.a(buffered_input), .b(12'b000111010111), .eq(weq471));
    equaln #(12) e472(.a(buffered_input), .b(12'b000111011000), .eq(weq472));
    equaln #(12) e473(.a(buffered_input), .b(12'b000111011001), .eq(weq473));
    equaln #(12) e474(.a(buffered_input), .b(12'b000111011010), .eq(weq474));
    equaln #(12) e475(.a(buffered_input), .b(12'b000111011011), .eq(weq475));
    equaln #(12) e476(.a(buffered_input), .b(12'b000111011100), .eq(weq476));
    equaln #(12) e477(.a(buffered_input), .b(12'b000111011101), .eq(weq477));
    equaln #(12) e478(.a(buffered_input), .b(12'b000111011110), .eq(weq478));
    equaln #(12) e479(.a(buffered_input), .b(12'b000111011111), .eq(weq479));
    equaln #(12) e480(.a(buffered_input), .b(12'b000111100000), .eq(weq480));
    equaln #(12) e481(.a(buffered_input), .b(12'b000111100001), .eq(weq481));
    equaln #(12) e482(.a(buffered_input), .b(12'b000111100010), .eq(weq482));
    equaln #(12) e483(.a(buffered_input), .b(12'b000111100011), .eq(weq483));
    equaln #(12) e484(.a(buffered_input), .b(12'b000111100100), .eq(weq484));
    equaln #(12) e485(.a(buffered_input), .b(12'b000111100101), .eq(weq485));
    equaln #(12) e486(.a(buffered_input), .b(12'b000111100110), .eq(weq486));
    equaln #(12) e487(.a(buffered_input), .b(12'b000111100111), .eq(weq487));
    equaln #(12) e488(.a(buffered_input), .b(12'b000111101000), .eq(weq488));
    equaln #(12) e489(.a(buffered_input), .b(12'b000111101001), .eq(weq489));
    equaln #(12) e490(.a(buffered_input), .b(12'b000111101010), .eq(weq490));
    equaln #(12) e491(.a(buffered_input), .b(12'b000111101011), .eq(weq491));
    equaln #(12) e492(.a(buffered_input), .b(12'b000111101100), .eq(weq492));
    equaln #(12) e493(.a(buffered_input), .b(12'b000111101101), .eq(weq493));
    equaln #(12) e494(.a(buffered_input), .b(12'b000111101110), .eq(weq494));
    equaln #(12) e495(.a(buffered_input), .b(12'b000111101111), .eq(weq495));
    equaln #(12) e496(.a(buffered_input), .b(12'b000111110000), .eq(weq496));
    equaln #(12) e497(.a(buffered_input), .b(12'b000111110001), .eq(weq497));
    equaln #(12) e498(.a(buffered_input), .b(12'b000111110010), .eq(weq498));
    equaln #(12) e499(.a(buffered_input), .b(12'b000111110011), .eq(weq499));
    equaln #(12) e500(.a(buffered_input), .b(12'b000111110100), .eq(weq500));
    equaln #(12) e501(.a(buffered_input), .b(12'b000111110101), .eq(weq501));
    equaln #(12) e502(.a(buffered_input), .b(12'b000111110110), .eq(weq502));
    equaln #(12) e503(.a(buffered_input), .b(12'b000111110111), .eq(weq503));
    equaln #(12) e504(.a(buffered_input), .b(12'b000111111000), .eq(weq504));
    equaln #(12) e505(.a(buffered_input), .b(12'b000111111001), .eq(weq505));
    equaln #(12) e506(.a(buffered_input), .b(12'b000111111010), .eq(weq506));
    equaln #(12) e507(.a(buffered_input), .b(12'b000111111011), .eq(weq507));
    equaln #(12) e508(.a(buffered_input), .b(12'b000111111100), .eq(weq508));
    equaln #(12) e509(.a(buffered_input), .b(12'b000111111101), .eq(weq509));
    equaln #(12) e510(.a(buffered_input), .b(12'b000111111110), .eq(weq510));
    equaln #(12) e511(.a(buffered_input), .b(12'b000111111111), .eq(weq511));
    equaln #(12) e512(.a(buffered_input), .b(12'b001000000000), .eq(weq512));
    equaln #(12) e513(.a(buffered_input), .b(12'b001000000001), .eq(weq513));
    equaln #(12) e514(.a(buffered_input), .b(12'b001000000010), .eq(weq514));
    equaln #(12) e515(.a(buffered_input), .b(12'b001000000011), .eq(weq515));
    equaln #(12) e516(.a(buffered_input), .b(12'b001000000100), .eq(weq516));
    equaln #(12) e517(.a(buffered_input), .b(12'b001000000101), .eq(weq517));
    equaln #(12) e518(.a(buffered_input), .b(12'b001000000110), .eq(weq518));
    equaln #(12) e519(.a(buffered_input), .b(12'b001000000111), .eq(weq519));
    equaln #(12) e520(.a(buffered_input), .b(12'b001000001000), .eq(weq520));
    equaln #(12) e521(.a(buffered_input), .b(12'b001000001001), .eq(weq521));
    equaln #(12) e522(.a(buffered_input), .b(12'b001000001010), .eq(weq522));
    equaln #(12) e523(.a(buffered_input), .b(12'b001000001011), .eq(weq523));
    equaln #(12) e524(.a(buffered_input), .b(12'b001000001100), .eq(weq524));
    equaln #(12) e525(.a(buffered_input), .b(12'b001000001101), .eq(weq525));
    equaln #(12) e526(.a(buffered_input), .b(12'b001000001110), .eq(weq526));
    equaln #(12) e527(.a(buffered_input), .b(12'b001000001111), .eq(weq527));
    equaln #(12) e528(.a(buffered_input), .b(12'b001000010000), .eq(weq528));
    equaln #(12) e529(.a(buffered_input), .b(12'b001000010001), .eq(weq529));
    equaln #(12) e530(.a(buffered_input), .b(12'b001000010010), .eq(weq530));
    equaln #(12) e531(.a(buffered_input), .b(12'b001000010011), .eq(weq531));
    equaln #(12) e532(.a(buffered_input), .b(12'b001000010100), .eq(weq532));
    equaln #(12) e533(.a(buffered_input), .b(12'b001000010101), .eq(weq533));
    equaln #(12) e534(.a(buffered_input), .b(12'b001000010110), .eq(weq534));
    equaln #(12) e535(.a(buffered_input), .b(12'b001000010111), .eq(weq535));
    equaln #(12) e536(.a(buffered_input), .b(12'b001000011000), .eq(weq536));
    equaln #(12) e537(.a(buffered_input), .b(12'b001000011001), .eq(weq537));
    equaln #(12) e538(.a(buffered_input), .b(12'b001000011010), .eq(weq538));
    equaln #(12) e539(.a(buffered_input), .b(12'b001000011011), .eq(weq539));
    equaln #(12) e540(.a(buffered_input), .b(12'b001000011100), .eq(weq540));
    equaln #(12) e541(.a(buffered_input), .b(12'b001000011101), .eq(weq541));
    equaln #(12) e542(.a(buffered_input), .b(12'b001000011110), .eq(weq542));
    equaln #(12) e543(.a(buffered_input), .b(12'b001000011111), .eq(weq543));
    equaln #(12) e544(.a(buffered_input), .b(12'b001000100000), .eq(weq544));
    equaln #(12) e545(.a(buffered_input), .b(12'b001000100001), .eq(weq545));
    equaln #(12) e546(.a(buffered_input), .b(12'b001000100010), .eq(weq546));
    equaln #(12) e547(.a(buffered_input), .b(12'b001000100011), .eq(weq547));
    equaln #(12) e548(.a(buffered_input), .b(12'b001000100100), .eq(weq548));
    equaln #(12) e549(.a(buffered_input), .b(12'b001000100101), .eq(weq549));
    equaln #(12) e550(.a(buffered_input), .b(12'b001000100110), .eq(weq550));
    equaln #(12) e551(.a(buffered_input), .b(12'b001000100111), .eq(weq551));
    equaln #(12) e552(.a(buffered_input), .b(12'b001000101000), .eq(weq552));
    equaln #(12) e553(.a(buffered_input), .b(12'b001000101001), .eq(weq553));
    equaln #(12) e554(.a(buffered_input), .b(12'b001000101010), .eq(weq554));
    equaln #(12) e555(.a(buffered_input), .b(12'b001000101011), .eq(weq555));
    equaln #(12) e556(.a(buffered_input), .b(12'b001000101100), .eq(weq556));
    equaln #(12) e557(.a(buffered_input), .b(12'b001000101101), .eq(weq557));
    equaln #(12) e558(.a(buffered_input), .b(12'b001000101110), .eq(weq558));
    equaln #(12) e559(.a(buffered_input), .b(12'b001000101111), .eq(weq559));
    equaln #(12) e560(.a(buffered_input), .b(12'b001000110000), .eq(weq560));
    equaln #(12) e561(.a(buffered_input), .b(12'b001000110001), .eq(weq561));
    equaln #(12) e562(.a(buffered_input), .b(12'b001000110010), .eq(weq562));
    equaln #(12) e563(.a(buffered_input), .b(12'b001000110011), .eq(weq563));
    equaln #(12) e564(.a(buffered_input), .b(12'b001000110100), .eq(weq564));
    equaln #(12) e565(.a(buffered_input), .b(12'b001000110101), .eq(weq565));
    equaln #(12) e566(.a(buffered_input), .b(12'b001000110110), .eq(weq566));
    equaln #(12) e567(.a(buffered_input), .b(12'b001000110111), .eq(weq567));
    equaln #(12) e568(.a(buffered_input), .b(12'b001000111000), .eq(weq568));
    equaln #(12) e569(.a(buffered_input), .b(12'b001000111001), .eq(weq569));
    equaln #(12) e570(.a(buffered_input), .b(12'b001000111010), .eq(weq570));
    equaln #(12) e571(.a(buffered_input), .b(12'b001000111011), .eq(weq571));
    equaln #(12) e572(.a(buffered_input), .b(12'b001000111100), .eq(weq572));
    equaln #(12) e573(.a(buffered_input), .b(12'b001000111101), .eq(weq573));
    equaln #(12) e574(.a(buffered_input), .b(12'b001000111110), .eq(weq574));
    equaln #(12) e575(.a(buffered_input), .b(12'b001000111111), .eq(weq575));
    equaln #(12) e576(.a(buffered_input), .b(12'b001001000000), .eq(weq576));
    equaln #(12) e577(.a(buffered_input), .b(12'b001001000001), .eq(weq577));
    equaln #(12) e578(.a(buffered_input), .b(12'b001001000010), .eq(weq578));
    equaln #(12) e579(.a(buffered_input), .b(12'b001001000011), .eq(weq579));
    equaln #(12) e580(.a(buffered_input), .b(12'b001001000100), .eq(weq580));
    equaln #(12) e581(.a(buffered_input), .b(12'b001001000101), .eq(weq581));
    equaln #(12) e582(.a(buffered_input), .b(12'b001001000110), .eq(weq582));
    equaln #(12) e583(.a(buffered_input), .b(12'b001001000111), .eq(weq583));
    equaln #(12) e584(.a(buffered_input), .b(12'b001001001000), .eq(weq584));
    equaln #(12) e585(.a(buffered_input), .b(12'b001001001001), .eq(weq585));
    equaln #(12) e586(.a(buffered_input), .b(12'b001001001010), .eq(weq586));
    equaln #(12) e587(.a(buffered_input), .b(12'b001001001011), .eq(weq587));
    equaln #(12) e588(.a(buffered_input), .b(12'b001001001100), .eq(weq588));
    equaln #(12) e589(.a(buffered_input), .b(12'b001001001101), .eq(weq589));
    equaln #(12) e590(.a(buffered_input), .b(12'b001001001110), .eq(weq590));
    equaln #(12) e591(.a(buffered_input), .b(12'b001001001111), .eq(weq591));
    equaln #(12) e592(.a(buffered_input), .b(12'b001001010000), .eq(weq592));
    equaln #(12) e593(.a(buffered_input), .b(12'b001001010001), .eq(weq593));
    equaln #(12) e594(.a(buffered_input), .b(12'b001001010010), .eq(weq594));
    equaln #(12) e595(.a(buffered_input), .b(12'b001001010011), .eq(weq595));
    equaln #(12) e596(.a(buffered_input), .b(12'b001001010100), .eq(weq596));
    equaln #(12) e597(.a(buffered_input), .b(12'b001001010101), .eq(weq597));
    equaln #(12) e598(.a(buffered_input), .b(12'b001001010110), .eq(weq598));
    equaln #(12) e599(.a(buffered_input), .b(12'b001001010111), .eq(weq599));
    equaln #(12) e600(.a(buffered_input), .b(12'b001001011000), .eq(weq600));
    equaln #(12) e601(.a(buffered_input), .b(12'b001001011001), .eq(weq601));
    equaln #(12) e602(.a(buffered_input), .b(12'b001001011010), .eq(weq602));
    equaln #(12) e603(.a(buffered_input), .b(12'b001001011011), .eq(weq603));
    equaln #(12) e604(.a(buffered_input), .b(12'b001001011100), .eq(weq604));
    equaln #(12) e605(.a(buffered_input), .b(12'b001001011101), .eq(weq605));
    equaln #(12) e606(.a(buffered_input), .b(12'b001001011110), .eq(weq606));
    equaln #(12) e607(.a(buffered_input), .b(12'b001001011111), .eq(weq607));
    equaln #(12) e608(.a(buffered_input), .b(12'b001001100000), .eq(weq608));
    equaln #(12) e609(.a(buffered_input), .b(12'b001001100001), .eq(weq609));
    equaln #(12) e610(.a(buffered_input), .b(12'b001001100010), .eq(weq610));
    equaln #(12) e611(.a(buffered_input), .b(12'b001001100011), .eq(weq611));
    equaln #(12) e612(.a(buffered_input), .b(12'b001001100100), .eq(weq612));
    equaln #(12) e613(.a(buffered_input), .b(12'b001001100101), .eq(weq613));
    equaln #(12) e614(.a(buffered_input), .b(12'b001001100110), .eq(weq614));
    equaln #(12) e615(.a(buffered_input), .b(12'b001001100111), .eq(weq615));
    equaln #(12) e616(.a(buffered_input), .b(12'b001001101000), .eq(weq616));
    equaln #(12) e617(.a(buffered_input), .b(12'b001001101001), .eq(weq617));
    equaln #(12) e618(.a(buffered_input), .b(12'b001001101010), .eq(weq618));
    equaln #(12) e619(.a(buffered_input), .b(12'b001001101011), .eq(weq619));
    equaln #(12) e620(.a(buffered_input), .b(12'b001001101100), .eq(weq620));
    equaln #(12) e621(.a(buffered_input), .b(12'b001001101101), .eq(weq621));
    equaln #(12) e622(.a(buffered_input), .b(12'b001001101110), .eq(weq622));
    equaln #(12) e623(.a(buffered_input), .b(12'b001001101111), .eq(weq623));
    equaln #(12) e624(.a(buffered_input), .b(12'b001001110000), .eq(weq624));
    equaln #(12) e625(.a(buffered_input), .b(12'b001001110001), .eq(weq625));
    equaln #(12) e626(.a(buffered_input), .b(12'b001001110010), .eq(weq626));
    equaln #(12) e627(.a(buffered_input), .b(12'b001001110011), .eq(weq627));
    equaln #(12) e628(.a(buffered_input), .b(12'b001001110100), .eq(weq628));
    equaln #(12) e629(.a(buffered_input), .b(12'b001001110101), .eq(weq629));
    equaln #(12) e630(.a(buffered_input), .b(12'b001001110110), .eq(weq630));
    equaln #(12) e631(.a(buffered_input), .b(12'b001001110111), .eq(weq631));
    equaln #(12) e632(.a(buffered_input), .b(12'b001001111000), .eq(weq632));
    equaln #(12) e633(.a(buffered_input), .b(12'b001001111001), .eq(weq633));
    equaln #(12) e634(.a(buffered_input), .b(12'b001001111010), .eq(weq634));
    equaln #(12) e635(.a(buffered_input), .b(12'b001001111011), .eq(weq635));
    equaln #(12) e636(.a(buffered_input), .b(12'b001001111100), .eq(weq636));
    equaln #(12) e637(.a(buffered_input), .b(12'b001001111101), .eq(weq637));
    equaln #(12) e638(.a(buffered_input), .b(12'b001001111110), .eq(weq638));
    equaln #(12) e639(.a(buffered_input), .b(12'b001001111111), .eq(weq639));
    equaln #(12) e640(.a(buffered_input), .b(12'b001010000000), .eq(weq640));
    equaln #(12) e641(.a(buffered_input), .b(12'b001010000001), .eq(weq641));
    equaln #(12) e642(.a(buffered_input), .b(12'b001010000010), .eq(weq642));
    equaln #(12) e643(.a(buffered_input), .b(12'b001010000011), .eq(weq643));
    equaln #(12) e644(.a(buffered_input), .b(12'b001010000100), .eq(weq644));
    equaln #(12) e645(.a(buffered_input), .b(12'b001010000101), .eq(weq645));
    equaln #(12) e646(.a(buffered_input), .b(12'b001010000110), .eq(weq646));
    equaln #(12) e647(.a(buffered_input), .b(12'b001010000111), .eq(weq647));
    equaln #(12) e648(.a(buffered_input), .b(12'b001010001000), .eq(weq648));
    equaln #(12) e649(.a(buffered_input), .b(12'b001010001001), .eq(weq649));
    equaln #(12) e650(.a(buffered_input), .b(12'b001010001010), .eq(weq650));
    equaln #(12) e651(.a(buffered_input), .b(12'b001010001011), .eq(weq651));
    equaln #(12) e652(.a(buffered_input), .b(12'b001010001100), .eq(weq652));
    equaln #(12) e653(.a(buffered_input), .b(12'b001010001101), .eq(weq653));
    equaln #(12) e654(.a(buffered_input), .b(12'b001010001110), .eq(weq654));
    equaln #(12) e655(.a(buffered_input), .b(12'b001010001111), .eq(weq655));
    equaln #(12) e656(.a(buffered_input), .b(12'b001010010000), .eq(weq656));
    equaln #(12) e657(.a(buffered_input), .b(12'b001010010001), .eq(weq657));
    equaln #(12) e658(.a(buffered_input), .b(12'b001010010010), .eq(weq658));
    equaln #(12) e659(.a(buffered_input), .b(12'b001010010011), .eq(weq659));
    equaln #(12) e660(.a(buffered_input), .b(12'b001010010100), .eq(weq660));
    equaln #(12) e661(.a(buffered_input), .b(12'b001010010101), .eq(weq661));
    equaln #(12) e662(.a(buffered_input), .b(12'b001010010110), .eq(weq662));
    equaln #(12) e663(.a(buffered_input), .b(12'b001010010111), .eq(weq663));
    equaln #(12) e664(.a(buffered_input), .b(12'b001010011000), .eq(weq664));
    equaln #(12) e665(.a(buffered_input), .b(12'b001010011001), .eq(weq665));
    equaln #(12) e666(.a(buffered_input), .b(12'b001010011010), .eq(weq666));
    equaln #(12) e667(.a(buffered_input), .b(12'b001010011011), .eq(weq667));
    equaln #(12) e668(.a(buffered_input), .b(12'b001010011100), .eq(weq668));
    equaln #(12) e669(.a(buffered_input), .b(12'b001010011101), .eq(weq669));
    equaln #(12) e670(.a(buffered_input), .b(12'b001010011110), .eq(weq670));
    equaln #(12) e671(.a(buffered_input), .b(12'b001010011111), .eq(weq671));
    equaln #(12) e672(.a(buffered_input), .b(12'b001010100000), .eq(weq672));
    equaln #(12) e673(.a(buffered_input), .b(12'b001010100001), .eq(weq673));
    equaln #(12) e674(.a(buffered_input), .b(12'b001010100010), .eq(weq674));
    equaln #(12) e675(.a(buffered_input), .b(12'b001010100011), .eq(weq675));
    equaln #(12) e676(.a(buffered_input), .b(12'b001010100100), .eq(weq676));
    equaln #(12) e677(.a(buffered_input), .b(12'b001010100101), .eq(weq677));
    equaln #(12) e678(.a(buffered_input), .b(12'b001010100110), .eq(weq678));
    equaln #(12) e679(.a(buffered_input), .b(12'b001010100111), .eq(weq679));
    equaln #(12) e680(.a(buffered_input), .b(12'b001010101000), .eq(weq680));
    equaln #(12) e681(.a(buffered_input), .b(12'b001010101001), .eq(weq681));
    equaln #(12) e682(.a(buffered_input), .b(12'b001010101010), .eq(weq682));
    equaln #(12) e683(.a(buffered_input), .b(12'b001010101011), .eq(weq683));
    equaln #(12) e684(.a(buffered_input), .b(12'b001010101100), .eq(weq684));
    equaln #(12) e685(.a(buffered_input), .b(12'b001010101101), .eq(weq685));
    equaln #(12) e686(.a(buffered_input), .b(12'b001010101110), .eq(weq686));
    equaln #(12) e687(.a(buffered_input), .b(12'b001010101111), .eq(weq687));
    equaln #(12) e688(.a(buffered_input), .b(12'b001010110000), .eq(weq688));
    equaln #(12) e689(.a(buffered_input), .b(12'b001010110001), .eq(weq689));
    equaln #(12) e690(.a(buffered_input), .b(12'b001010110010), .eq(weq690));
    equaln #(12) e691(.a(buffered_input), .b(12'b001010110011), .eq(weq691));
    equaln #(12) e692(.a(buffered_input), .b(12'b001010110100), .eq(weq692));
    equaln #(12) e693(.a(buffered_input), .b(12'b001010110101), .eq(weq693));
    equaln #(12) e694(.a(buffered_input), .b(12'b001010110110), .eq(weq694));
    equaln #(12) e695(.a(buffered_input), .b(12'b001010110111), .eq(weq695));
    equaln #(12) e696(.a(buffered_input), .b(12'b001010111000), .eq(weq696));
    equaln #(12) e697(.a(buffered_input), .b(12'b001010111001), .eq(weq697));
    equaln #(12) e698(.a(buffered_input), .b(12'b001010111010), .eq(weq698));
    equaln #(12) e699(.a(buffered_input), .b(12'b001010111011), .eq(weq699));
    equaln #(12) e700(.a(buffered_input), .b(12'b001010111100), .eq(weq700));
    equaln #(12) e701(.a(buffered_input), .b(12'b001010111101), .eq(weq701));
    equaln #(12) e702(.a(buffered_input), .b(12'b001010111110), .eq(weq702));
    equaln #(12) e703(.a(buffered_input), .b(12'b001010111111), .eq(weq703));
    equaln #(12) e704(.a(buffered_input), .b(12'b001011000000), .eq(weq704));
    equaln #(12) e705(.a(buffered_input), .b(12'b001011000001), .eq(weq705));
    equaln #(12) e706(.a(buffered_input), .b(12'b001011000010), .eq(weq706));
    equaln #(12) e707(.a(buffered_input), .b(12'b001011000011), .eq(weq707));
    equaln #(12) e708(.a(buffered_input), .b(12'b001011000100), .eq(weq708));
    equaln #(12) e709(.a(buffered_input), .b(12'b001011000101), .eq(weq709));
    equaln #(12) e710(.a(buffered_input), .b(12'b001011000110), .eq(weq710));
    equaln #(12) e711(.a(buffered_input), .b(12'b001011000111), .eq(weq711));
    equaln #(12) e712(.a(buffered_input), .b(12'b001011001000), .eq(weq712));
    equaln #(12) e713(.a(buffered_input), .b(12'b001011001001), .eq(weq713));
    equaln #(12) e714(.a(buffered_input), .b(12'b001011001010), .eq(weq714));
    equaln #(12) e715(.a(buffered_input), .b(12'b001011001011), .eq(weq715));
    equaln #(12) e716(.a(buffered_input), .b(12'b001011001100), .eq(weq716));
    equaln #(12) e717(.a(buffered_input), .b(12'b001011001101), .eq(weq717));
    equaln #(12) e718(.a(buffered_input), .b(12'b001011001110), .eq(weq718));
    equaln #(12) e719(.a(buffered_input), .b(12'b001011001111), .eq(weq719));
    equaln #(12) e720(.a(buffered_input), .b(12'b001011010000), .eq(weq720));
    equaln #(12) e721(.a(buffered_input), .b(12'b001011010001), .eq(weq721));
    equaln #(12) e722(.a(buffered_input), .b(12'b001011010010), .eq(weq722));
    equaln #(12) e723(.a(buffered_input), .b(12'b001011010011), .eq(weq723));
    equaln #(12) e724(.a(buffered_input), .b(12'b001011010100), .eq(weq724));
    equaln #(12) e725(.a(buffered_input), .b(12'b001011010101), .eq(weq725));
    equaln #(12) e726(.a(buffered_input), .b(12'b001011010110), .eq(weq726));
    equaln #(12) e727(.a(buffered_input), .b(12'b001011010111), .eq(weq727));
    equaln #(12) e728(.a(buffered_input), .b(12'b001011011000), .eq(weq728));
    equaln #(12) e729(.a(buffered_input), .b(12'b001011011001), .eq(weq729));
    equaln #(12) e730(.a(buffered_input), .b(12'b001011011010), .eq(weq730));
    equaln #(12) e731(.a(buffered_input), .b(12'b001011011011), .eq(weq731));
    equaln #(12) e732(.a(buffered_input), .b(12'b001011011100), .eq(weq732));
    equaln #(12) e733(.a(buffered_input), .b(12'b001011011101), .eq(weq733));
    equaln #(12) e734(.a(buffered_input), .b(12'b001011011110), .eq(weq734));
    equaln #(12) e735(.a(buffered_input), .b(12'b001011011111), .eq(weq735));
    equaln #(12) e736(.a(buffered_input), .b(12'b001011100000), .eq(weq736));
    equaln #(12) e737(.a(buffered_input), .b(12'b001011100001), .eq(weq737));
    equaln #(12) e738(.a(buffered_input), .b(12'b001011100010), .eq(weq738));
    equaln #(12) e739(.a(buffered_input), .b(12'b001011100011), .eq(weq739));
    equaln #(12) e740(.a(buffered_input), .b(12'b001011100100), .eq(weq740));
    equaln #(12) e741(.a(buffered_input), .b(12'b001011100101), .eq(weq741));
    equaln #(12) e742(.a(buffered_input), .b(12'b001011100110), .eq(weq742));
    equaln #(12) e743(.a(buffered_input), .b(12'b001011100111), .eq(weq743));
    equaln #(12) e744(.a(buffered_input), .b(12'b001011101000), .eq(weq744));
    equaln #(12) e745(.a(buffered_input), .b(12'b001011101001), .eq(weq745));
    equaln #(12) e746(.a(buffered_input), .b(12'b001011101010), .eq(weq746));
    equaln #(12) e747(.a(buffered_input), .b(12'b001011101011), .eq(weq747));
    equaln #(12) e748(.a(buffered_input), .b(12'b001011101100), .eq(weq748));
    equaln #(12) e749(.a(buffered_input), .b(12'b001011101101), .eq(weq749));
    equaln #(12) e750(.a(buffered_input), .b(12'b001011101110), .eq(weq750));
    equaln #(12) e751(.a(buffered_input), .b(12'b001011101111), .eq(weq751));
    equaln #(12) e752(.a(buffered_input), .b(12'b001011110000), .eq(weq752));
    equaln #(12) e753(.a(buffered_input), .b(12'b001011110001), .eq(weq753));
    equaln #(12) e754(.a(buffered_input), .b(12'b001011110010), .eq(weq754));
    equaln #(12) e755(.a(buffered_input), .b(12'b001011110011), .eq(weq755));
    equaln #(12) e756(.a(buffered_input), .b(12'b001011110100), .eq(weq756));
    equaln #(12) e757(.a(buffered_input), .b(12'b001011110101), .eq(weq757));
    equaln #(12) e758(.a(buffered_input), .b(12'b001011110110), .eq(weq758));
    equaln #(12) e759(.a(buffered_input), .b(12'b001011110111), .eq(weq759));
    equaln #(12) e760(.a(buffered_input), .b(12'b001011111000), .eq(weq760));
    equaln #(12) e761(.a(buffered_input), .b(12'b001011111001), .eq(weq761));
    equaln #(12) e762(.a(buffered_input), .b(12'b001011111010), .eq(weq762));
    equaln #(12) e763(.a(buffered_input), .b(12'b001011111011), .eq(weq763));
    equaln #(12) e764(.a(buffered_input), .b(12'b001011111100), .eq(weq764));
    equaln #(12) e765(.a(buffered_input), .b(12'b001011111101), .eq(weq765));
    equaln #(12) e766(.a(buffered_input), .b(12'b001011111110), .eq(weq766));
    equaln #(12) e767(.a(buffered_input), .b(12'b001011111111), .eq(weq767));
    equaln #(12) e768(.a(buffered_input), .b(12'b001100000000), .eq(weq768));
    equaln #(12) e769(.a(buffered_input), .b(12'b001100000001), .eq(weq769));
    equaln #(12) e770(.a(buffered_input), .b(12'b001100000010), .eq(weq770));
    equaln #(12) e771(.a(buffered_input), .b(12'b001100000011), .eq(weq771));
    equaln #(12) e772(.a(buffered_input), .b(12'b001100000100), .eq(weq772));
    equaln #(12) e773(.a(buffered_input), .b(12'b001100000101), .eq(weq773));
    equaln #(12) e774(.a(buffered_input), .b(12'b001100000110), .eq(weq774));
    equaln #(12) e775(.a(buffered_input), .b(12'b001100000111), .eq(weq775));
    equaln #(12) e776(.a(buffered_input), .b(12'b001100001000), .eq(weq776));
    equaln #(12) e777(.a(buffered_input), .b(12'b001100001001), .eq(weq777));
    equaln #(12) e778(.a(buffered_input), .b(12'b001100001010), .eq(weq778));
    equaln #(12) e779(.a(buffered_input), .b(12'b001100001011), .eq(weq779));
    equaln #(12) e780(.a(buffered_input), .b(12'b001100001100), .eq(weq780));
    equaln #(12) e781(.a(buffered_input), .b(12'b001100001101), .eq(weq781));
    equaln #(12) e782(.a(buffered_input), .b(12'b001100001110), .eq(weq782));
    equaln #(12) e783(.a(buffered_input), .b(12'b001100001111), .eq(weq783));
    equaln #(12) e784(.a(buffered_input), .b(12'b001100010000), .eq(weq784));
    equaln #(12) e785(.a(buffered_input), .b(12'b001100010001), .eq(weq785));
    equaln #(12) e786(.a(buffered_input), .b(12'b001100010010), .eq(weq786));
    equaln #(12) e787(.a(buffered_input), .b(12'b001100010011), .eq(weq787));
    equaln #(12) e788(.a(buffered_input), .b(12'b001100010100), .eq(weq788));
    equaln #(12) e789(.a(buffered_input), .b(12'b001100010101), .eq(weq789));
    equaln #(12) e790(.a(buffered_input), .b(12'b001100010110), .eq(weq790));
    equaln #(12) e791(.a(buffered_input), .b(12'b001100010111), .eq(weq791));
    equaln #(12) e792(.a(buffered_input), .b(12'b001100011000), .eq(weq792));
    equaln #(12) e793(.a(buffered_input), .b(12'b001100011001), .eq(weq793));
    equaln #(12) e794(.a(buffered_input), .b(12'b001100011010), .eq(weq794));
    equaln #(12) e795(.a(buffered_input), .b(12'b001100011011), .eq(weq795));
    equaln #(12) e796(.a(buffered_input), .b(12'b001100011100), .eq(weq796));
    equaln #(12) e797(.a(buffered_input), .b(12'b001100011101), .eq(weq797));
    equaln #(12) e798(.a(buffered_input), .b(12'b001100011110), .eq(weq798));
    equaln #(12) e799(.a(buffered_input), .b(12'b001100011111), .eq(weq799));
    equaln #(12) e800(.a(buffered_input), .b(12'b001100100000), .eq(weq800));
    equaln #(12) e801(.a(buffered_input), .b(12'b001100100001), .eq(weq801));
    equaln #(12) e802(.a(buffered_input), .b(12'b001100100010), .eq(weq802));
    equaln #(12) e803(.a(buffered_input), .b(12'b001100100011), .eq(weq803));
    equaln #(12) e804(.a(buffered_input), .b(12'b001100100100), .eq(weq804));
    equaln #(12) e805(.a(buffered_input), .b(12'b001100100101), .eq(weq805));
    equaln #(12) e806(.a(buffered_input), .b(12'b001100100110), .eq(weq806));
    equaln #(12) e807(.a(buffered_input), .b(12'b001100100111), .eq(weq807));
    equaln #(12) e808(.a(buffered_input), .b(12'b001100101000), .eq(weq808));
    equaln #(12) e809(.a(buffered_input), .b(12'b001100101001), .eq(weq809));
    equaln #(12) e810(.a(buffered_input), .b(12'b001100101010), .eq(weq810));
    equaln #(12) e811(.a(buffered_input), .b(12'b001100101011), .eq(weq811));
    equaln #(12) e812(.a(buffered_input), .b(12'b001100101100), .eq(weq812));
    equaln #(12) e813(.a(buffered_input), .b(12'b001100101101), .eq(weq813));
    equaln #(12) e814(.a(buffered_input), .b(12'b001100101110), .eq(weq814));
    equaln #(12) e815(.a(buffered_input), .b(12'b001100101111), .eq(weq815));
    equaln #(12) e816(.a(buffered_input), .b(12'b001100110000), .eq(weq816));
    equaln #(12) e817(.a(buffered_input), .b(12'b001100110001), .eq(weq817));
    equaln #(12) e818(.a(buffered_input), .b(12'b001100110010), .eq(weq818));
    equaln #(12) e819(.a(buffered_input), .b(12'b001100110011), .eq(weq819));
    equaln #(12) e820(.a(buffered_input), .b(12'b001100110100), .eq(weq820));
    equaln #(12) e821(.a(buffered_input), .b(12'b001100110101), .eq(weq821));
    equaln #(12) e822(.a(buffered_input), .b(12'b001100110110), .eq(weq822));
    equaln #(12) e823(.a(buffered_input), .b(12'b001100110111), .eq(weq823));
    equaln #(12) e824(.a(buffered_input), .b(12'b001100111000), .eq(weq824));
    equaln #(12) e825(.a(buffered_input), .b(12'b001100111001), .eq(weq825));
    equaln #(12) e826(.a(buffered_input), .b(12'b001100111010), .eq(weq826));
    equaln #(12) e827(.a(buffered_input), .b(12'b001100111011), .eq(weq827));
    equaln #(12) e828(.a(buffered_input), .b(12'b001100111100), .eq(weq828));
    equaln #(12) e829(.a(buffered_input), .b(12'b001100111101), .eq(weq829));
    equaln #(12) e830(.a(buffered_input), .b(12'b001100111110), .eq(weq830));
    equaln #(12) e831(.a(buffered_input), .b(12'b001100111111), .eq(weq831));
    equaln #(12) e832(.a(buffered_input), .b(12'b001101000000), .eq(weq832));
    equaln #(12) e833(.a(buffered_input), .b(12'b001101000001), .eq(weq833));
    equaln #(12) e834(.a(buffered_input), .b(12'b001101000010), .eq(weq834));
    equaln #(12) e835(.a(buffered_input), .b(12'b001101000011), .eq(weq835));
    equaln #(12) e836(.a(buffered_input), .b(12'b001101000100), .eq(weq836));
    equaln #(12) e837(.a(buffered_input), .b(12'b001101000101), .eq(weq837));
    equaln #(12) e838(.a(buffered_input), .b(12'b001101000110), .eq(weq838));
    equaln #(12) e839(.a(buffered_input), .b(12'b001101000111), .eq(weq839));
    equaln #(12) e840(.a(buffered_input), .b(12'b001101001000), .eq(weq840));
    equaln #(12) e841(.a(buffered_input), .b(12'b001101001001), .eq(weq841));
    equaln #(12) e842(.a(buffered_input), .b(12'b001101001010), .eq(weq842));
    equaln #(12) e843(.a(buffered_input), .b(12'b001101001011), .eq(weq843));
    equaln #(12) e844(.a(buffered_input), .b(12'b001101001100), .eq(weq844));
    equaln #(12) e845(.a(buffered_input), .b(12'b001101001101), .eq(weq845));
    equaln #(12) e846(.a(buffered_input), .b(12'b001101001110), .eq(weq846));
    equaln #(12) e847(.a(buffered_input), .b(12'b001101001111), .eq(weq847));
    equaln #(12) e848(.a(buffered_input), .b(12'b001101010000), .eq(weq848));
    equaln #(12) e849(.a(buffered_input), .b(12'b001101010001), .eq(weq849));
    equaln #(12) e850(.a(buffered_input), .b(12'b001101010010), .eq(weq850));
    equaln #(12) e851(.a(buffered_input), .b(12'b001101010011), .eq(weq851));
    equaln #(12) e852(.a(buffered_input), .b(12'b001101010100), .eq(weq852));
    equaln #(12) e853(.a(buffered_input), .b(12'b001101010101), .eq(weq853));
    equaln #(12) e854(.a(buffered_input), .b(12'b001101010110), .eq(weq854));
    equaln #(12) e855(.a(buffered_input), .b(12'b001101010111), .eq(weq855));
    equaln #(12) e856(.a(buffered_input), .b(12'b001101011000), .eq(weq856));
    equaln #(12) e857(.a(buffered_input), .b(12'b001101011001), .eq(weq857));
    equaln #(12) e858(.a(buffered_input), .b(12'b001101011010), .eq(weq858));
    equaln #(12) e859(.a(buffered_input), .b(12'b001101011011), .eq(weq859));
    equaln #(12) e860(.a(buffered_input), .b(12'b001101011100), .eq(weq860));
    equaln #(12) e861(.a(buffered_input), .b(12'b001101011101), .eq(weq861));
    equaln #(12) e862(.a(buffered_input), .b(12'b001101011110), .eq(weq862));
    equaln #(12) e863(.a(buffered_input), .b(12'b001101011111), .eq(weq863));
    equaln #(12) e864(.a(buffered_input), .b(12'b001101100000), .eq(weq864));
    equaln #(12) e865(.a(buffered_input), .b(12'b001101100001), .eq(weq865));
    equaln #(12) e866(.a(buffered_input), .b(12'b001101100010), .eq(weq866));
    equaln #(12) e867(.a(buffered_input), .b(12'b001101100011), .eq(weq867));
    equaln #(12) e868(.a(buffered_input), .b(12'b001101100100), .eq(weq868));
    equaln #(12) e869(.a(buffered_input), .b(12'b001101100101), .eq(weq869));
    equaln #(12) e870(.a(buffered_input), .b(12'b001101100110), .eq(weq870));
    equaln #(12) e871(.a(buffered_input), .b(12'b001101100111), .eq(weq871));
    equaln #(12) e872(.a(buffered_input), .b(12'b001101101000), .eq(weq872));
    equaln #(12) e873(.a(buffered_input), .b(12'b001101101001), .eq(weq873));
    equaln #(12) e874(.a(buffered_input), .b(12'b001101101010), .eq(weq874));
    equaln #(12) e875(.a(buffered_input), .b(12'b001101101011), .eq(weq875));
    equaln #(12) e876(.a(buffered_input), .b(12'b001101101100), .eq(weq876));
    equaln #(12) e877(.a(buffered_input), .b(12'b001101101101), .eq(weq877));
    equaln #(12) e878(.a(buffered_input), .b(12'b001101101110), .eq(weq878));
    equaln #(12) e879(.a(buffered_input), .b(12'b001101101111), .eq(weq879));
    equaln #(12) e880(.a(buffered_input), .b(12'b001101110000), .eq(weq880));
    equaln #(12) e881(.a(buffered_input), .b(12'b001101110001), .eq(weq881));
    equaln #(12) e882(.a(buffered_input), .b(12'b001101110010), .eq(weq882));
    equaln #(12) e883(.a(buffered_input), .b(12'b001101110011), .eq(weq883));
    equaln #(12) e884(.a(buffered_input), .b(12'b001101110100), .eq(weq884));
    equaln #(12) e885(.a(buffered_input), .b(12'b001101110101), .eq(weq885));
    equaln #(12) e886(.a(buffered_input), .b(12'b001101110110), .eq(weq886));
    equaln #(12) e887(.a(buffered_input), .b(12'b001101110111), .eq(weq887));
    equaln #(12) e888(.a(buffered_input), .b(12'b001101111000), .eq(weq888));
    equaln #(12) e889(.a(buffered_input), .b(12'b001101111001), .eq(weq889));
    equaln #(12) e890(.a(buffered_input), .b(12'b001101111010), .eq(weq890));
    equaln #(12) e891(.a(buffered_input), .b(12'b001101111011), .eq(weq891));
    equaln #(12) e892(.a(buffered_input), .b(12'b001101111100), .eq(weq892));
    equaln #(12) e893(.a(buffered_input), .b(12'b001101111101), .eq(weq893));
    equaln #(12) e894(.a(buffered_input), .b(12'b001101111110), .eq(weq894));
    equaln #(12) e895(.a(buffered_input), .b(12'b001101111111), .eq(weq895));
    equaln #(12) e896(.a(buffered_input), .b(12'b001110000000), .eq(weq896));
    equaln #(12) e897(.a(buffered_input), .b(12'b001110000001), .eq(weq897));
    equaln #(12) e898(.a(buffered_input), .b(12'b001110000010), .eq(weq898));
    equaln #(12) e899(.a(buffered_input), .b(12'b001110000011), .eq(weq899));
    equaln #(12) e900(.a(buffered_input), .b(12'b001110000100), .eq(weq900));
    equaln #(12) e901(.a(buffered_input), .b(12'b001110000101), .eq(weq901));
    equaln #(12) e902(.a(buffered_input), .b(12'b001110000110), .eq(weq902));
    equaln #(12) e903(.a(buffered_input), .b(12'b001110000111), .eq(weq903));
    equaln #(12) e904(.a(buffered_input), .b(12'b001110001000), .eq(weq904));
    equaln #(12) e905(.a(buffered_input), .b(12'b001110001001), .eq(weq905));
    equaln #(12) e906(.a(buffered_input), .b(12'b001110001010), .eq(weq906));
    equaln #(12) e907(.a(buffered_input), .b(12'b001110001011), .eq(weq907));
    equaln #(12) e908(.a(buffered_input), .b(12'b001110001100), .eq(weq908));
    equaln #(12) e909(.a(buffered_input), .b(12'b001110001101), .eq(weq909));
    equaln #(12) e910(.a(buffered_input), .b(12'b001110001110), .eq(weq910));
    equaln #(12) e911(.a(buffered_input), .b(12'b001110001111), .eq(weq911));
    equaln #(12) e912(.a(buffered_input), .b(12'b001110010000), .eq(weq912));
    equaln #(12) e913(.a(buffered_input), .b(12'b001110010001), .eq(weq913));
    equaln #(12) e914(.a(buffered_input), .b(12'b001110010010), .eq(weq914));
    equaln #(12) e915(.a(buffered_input), .b(12'b001110010011), .eq(weq915));
    equaln #(12) e916(.a(buffered_input), .b(12'b001110010100), .eq(weq916));
    equaln #(12) e917(.a(buffered_input), .b(12'b001110010101), .eq(weq917));
    equaln #(12) e918(.a(buffered_input), .b(12'b001110010110), .eq(weq918));
    equaln #(12) e919(.a(buffered_input), .b(12'b001110010111), .eq(weq919));
    equaln #(12) e920(.a(buffered_input), .b(12'b001110011000), .eq(weq920));
    equaln #(12) e921(.a(buffered_input), .b(12'b001110011001), .eq(weq921));
    equaln #(12) e922(.a(buffered_input), .b(12'b001110011010), .eq(weq922));
    equaln #(12) e923(.a(buffered_input), .b(12'b001110011011), .eq(weq923));
    equaln #(12) e924(.a(buffered_input), .b(12'b001110011100), .eq(weq924));
    equaln #(12) e925(.a(buffered_input), .b(12'b001110011101), .eq(weq925));
    equaln #(12) e926(.a(buffered_input), .b(12'b001110011110), .eq(weq926));
    equaln #(12) e927(.a(buffered_input), .b(12'b001110011111), .eq(weq927));
    equaln #(12) e928(.a(buffered_input), .b(12'b001110100000), .eq(weq928));
    equaln #(12) e929(.a(buffered_input), .b(12'b001110100001), .eq(weq929));
    equaln #(12) e930(.a(buffered_input), .b(12'b001110100010), .eq(weq930));
    equaln #(12) e931(.a(buffered_input), .b(12'b001110100011), .eq(weq931));
    equaln #(12) e932(.a(buffered_input), .b(12'b001110100100), .eq(weq932));
    equaln #(12) e933(.a(buffered_input), .b(12'b001110100101), .eq(weq933));
    equaln #(12) e934(.a(buffered_input), .b(12'b001110100110), .eq(weq934));
    equaln #(12) e935(.a(buffered_input), .b(12'b001110100111), .eq(weq935));
    equaln #(12) e936(.a(buffered_input), .b(12'b001110101000), .eq(weq936));
    equaln #(12) e937(.a(buffered_input), .b(12'b001110101001), .eq(weq937));
    equaln #(12) e938(.a(buffered_input), .b(12'b001110101010), .eq(weq938));
    equaln #(12) e939(.a(buffered_input), .b(12'b001110101011), .eq(weq939));
    equaln #(12) e940(.a(buffered_input), .b(12'b001110101100), .eq(weq940));
    equaln #(12) e941(.a(buffered_input), .b(12'b001110101101), .eq(weq941));
    equaln #(12) e942(.a(buffered_input), .b(12'b001110101110), .eq(weq942));
    equaln #(12) e943(.a(buffered_input), .b(12'b001110101111), .eq(weq943));
    equaln #(12) e944(.a(buffered_input), .b(12'b001110110000), .eq(weq944));
    equaln #(12) e945(.a(buffered_input), .b(12'b001110110001), .eq(weq945));
    equaln #(12) e946(.a(buffered_input), .b(12'b001110110010), .eq(weq946));
    equaln #(12) e947(.a(buffered_input), .b(12'b001110110011), .eq(weq947));
    equaln #(12) e948(.a(buffered_input), .b(12'b001110110100), .eq(weq948));
    equaln #(12) e949(.a(buffered_input), .b(12'b001110110101), .eq(weq949));
    equaln #(12) e950(.a(buffered_input), .b(12'b001110110110), .eq(weq950));
    equaln #(12) e951(.a(buffered_input), .b(12'b001110110111), .eq(weq951));
    equaln #(12) e952(.a(buffered_input), .b(12'b001110111000), .eq(weq952));
    equaln #(12) e953(.a(buffered_input), .b(12'b001110111001), .eq(weq953));
    equaln #(12) e954(.a(buffered_input), .b(12'b001110111010), .eq(weq954));
    equaln #(12) e955(.a(buffered_input), .b(12'b001110111011), .eq(weq955));
    equaln #(12) e956(.a(buffered_input), .b(12'b001110111100), .eq(weq956));
    equaln #(12) e957(.a(buffered_input), .b(12'b001110111101), .eq(weq957));
    equaln #(12) e958(.a(buffered_input), .b(12'b001110111110), .eq(weq958));
    equaln #(12) e959(.a(buffered_input), .b(12'b001110111111), .eq(weq959));
    equaln #(12) e960(.a(buffered_input), .b(12'b001111000000), .eq(weq960));
    equaln #(12) e961(.a(buffered_input), .b(12'b001111000001), .eq(weq961));
    equaln #(12) e962(.a(buffered_input), .b(12'b001111000010), .eq(weq962));
    equaln #(12) e963(.a(buffered_input), .b(12'b001111000011), .eq(weq963));
    equaln #(12) e964(.a(buffered_input), .b(12'b001111000100), .eq(weq964));
    equaln #(12) e965(.a(buffered_input), .b(12'b001111000101), .eq(weq965));
    equaln #(12) e966(.a(buffered_input), .b(12'b001111000110), .eq(weq966));
    equaln #(12) e967(.a(buffered_input), .b(12'b001111000111), .eq(weq967));
    equaln #(12) e968(.a(buffered_input), .b(12'b001111001000), .eq(weq968));
    equaln #(12) e969(.a(buffered_input), .b(12'b001111001001), .eq(weq969));
    equaln #(12) e970(.a(buffered_input), .b(12'b001111001010), .eq(weq970));
    equaln #(12) e971(.a(buffered_input), .b(12'b001111001011), .eq(weq971));
    equaln #(12) e972(.a(buffered_input), .b(12'b001111001100), .eq(weq972));
    equaln #(12) e973(.a(buffered_input), .b(12'b001111001101), .eq(weq973));
    equaln #(12) e974(.a(buffered_input), .b(12'b001111001110), .eq(weq974));
    equaln #(12) e975(.a(buffered_input), .b(12'b001111001111), .eq(weq975));
    equaln #(12) e976(.a(buffered_input), .b(12'b001111010000), .eq(weq976));
    equaln #(12) e977(.a(buffered_input), .b(12'b001111010001), .eq(weq977));
    equaln #(12) e978(.a(buffered_input), .b(12'b001111010010), .eq(weq978));
    equaln #(12) e979(.a(buffered_input), .b(12'b001111010011), .eq(weq979));
    equaln #(12) e980(.a(buffered_input), .b(12'b001111010100), .eq(weq980));
    equaln #(12) e981(.a(buffered_input), .b(12'b001111010101), .eq(weq981));
    equaln #(12) e982(.a(buffered_input), .b(12'b001111010110), .eq(weq982));
    equaln #(12) e983(.a(buffered_input), .b(12'b001111010111), .eq(weq983));
    equaln #(12) e984(.a(buffered_input), .b(12'b001111011000), .eq(weq984));
    equaln #(12) e985(.a(buffered_input), .b(12'b001111011001), .eq(weq985));
    equaln #(12) e986(.a(buffered_input), .b(12'b001111011010), .eq(weq986));
    equaln #(12) e987(.a(buffered_input), .b(12'b001111011011), .eq(weq987));
    equaln #(12) e988(.a(buffered_input), .b(12'b001111011100), .eq(weq988));
    equaln #(12) e989(.a(buffered_input), .b(12'b001111011101), .eq(weq989));
    equaln #(12) e990(.a(buffered_input), .b(12'b001111011110), .eq(weq990));
    equaln #(12) e991(.a(buffered_input), .b(12'b001111011111), .eq(weq991));
    equaln #(12) e992(.a(buffered_input), .b(12'b001111100000), .eq(weq992));
    equaln #(12) e993(.a(buffered_input), .b(12'b001111100001), .eq(weq993));
    equaln #(12) e994(.a(buffered_input), .b(12'b001111100010), .eq(weq994));
    equaln #(12) e995(.a(buffered_input), .b(12'b001111100011), .eq(weq995));
    equaln #(12) e996(.a(buffered_input), .b(12'b001111100100), .eq(weq996));
    equaln #(12) e997(.a(buffered_input), .b(12'b001111100101), .eq(weq997));
    equaln #(12) e998(.a(buffered_input), .b(12'b001111100110), .eq(weq998));
    equaln #(12) e999(.a(buffered_input), .b(12'b001111100111), .eq(weq999));
    equaln #(12) e1000(.a(buffered_input), .b(12'b001111101000), .eq(weq1000));
    equaln #(12) e1001(.a(buffered_input), .b(12'b001111101001), .eq(weq1001));
    equaln #(12) e1002(.a(buffered_input), .b(12'b001111101010), .eq(weq1002));
    equaln #(12) e1003(.a(buffered_input), .b(12'b001111101011), .eq(weq1003));
    equaln #(12) e1004(.a(buffered_input), .b(12'b001111101100), .eq(weq1004));
    equaln #(12) e1005(.a(buffered_input), .b(12'b001111101101), .eq(weq1005));
    equaln #(12) e1006(.a(buffered_input), .b(12'b001111101110), .eq(weq1006));
    equaln #(12) e1007(.a(buffered_input), .b(12'b001111101111), .eq(weq1007));
    equaln #(12) e1008(.a(buffered_input), .b(12'b001111110000), .eq(weq1008));
    equaln #(12) e1009(.a(buffered_input), .b(12'b001111110001), .eq(weq1009));
    equaln #(12) e1010(.a(buffered_input), .b(12'b001111110010), .eq(weq1010));
    equaln #(12) e1011(.a(buffered_input), .b(12'b001111110011), .eq(weq1011));
    equaln #(12) e1012(.a(buffered_input), .b(12'b001111110100), .eq(weq1012));
    equaln #(12) e1013(.a(buffered_input), .b(12'b001111110101), .eq(weq1013));
    equaln #(12) e1014(.a(buffered_input), .b(12'b001111110110), .eq(weq1014));
    equaln #(12) e1015(.a(buffered_input), .b(12'b001111110111), .eq(weq1015));
    equaln #(12) e1016(.a(buffered_input), .b(12'b001111111000), .eq(weq1016));
    equaln #(12) e1017(.a(buffered_input), .b(12'b001111111001), .eq(weq1017));
    equaln #(12) e1018(.a(buffered_input), .b(12'b001111111010), .eq(weq1018));
    equaln #(12) e1019(.a(buffered_input), .b(12'b001111111011), .eq(weq1019));
    equaln #(12) e1020(.a(buffered_input), .b(12'b001111111100), .eq(weq1020));
    equaln #(12) e1021(.a(buffered_input), .b(12'b001111111101), .eq(weq1021));
    equaln #(12) e1022(.a(buffered_input), .b(12'b001111111110), .eq(weq1022));
    equaln #(12) e1023(.a(buffered_input), .b(12'b001111111111), .eq(weq1023));
    equaln #(12) e1024(.a(buffered_input), .b(12'b010000000000), .eq(weq1024));
    equaln #(12) e1025(.a(buffered_input), .b(12'b010000000001), .eq(weq1025));
    equaln #(12) e1026(.a(buffered_input), .b(12'b010000000010), .eq(weq1026));
    equaln #(12) e1027(.a(buffered_input), .b(12'b010000000011), .eq(weq1027));
    equaln #(12) e1028(.a(buffered_input), .b(12'b010000000100), .eq(weq1028));
    equaln #(12) e1029(.a(buffered_input), .b(12'b010000000101), .eq(weq1029));
    equaln #(12) e1030(.a(buffered_input), .b(12'b010000000110), .eq(weq1030));
    equaln #(12) e1031(.a(buffered_input), .b(12'b010000000111), .eq(weq1031));
    equaln #(12) e1032(.a(buffered_input), .b(12'b010000001000), .eq(weq1032));
    equaln #(12) e1033(.a(buffered_input), .b(12'b010000001001), .eq(weq1033));
    equaln #(12) e1034(.a(buffered_input), .b(12'b010000001010), .eq(weq1034));
    equaln #(12) e1035(.a(buffered_input), .b(12'b010000001011), .eq(weq1035));
    equaln #(12) e1036(.a(buffered_input), .b(12'b010000001100), .eq(weq1036));
    equaln #(12) e1037(.a(buffered_input), .b(12'b010000001101), .eq(weq1037));
    equaln #(12) e1038(.a(buffered_input), .b(12'b010000001110), .eq(weq1038));
    equaln #(12) e1039(.a(buffered_input), .b(12'b010000001111), .eq(weq1039));
    equaln #(12) e1040(.a(buffered_input), .b(12'b010000010000), .eq(weq1040));
    equaln #(12) e1041(.a(buffered_input), .b(12'b010000010001), .eq(weq1041));
    equaln #(12) e1042(.a(buffered_input), .b(12'b010000010010), .eq(weq1042));
    equaln #(12) e1043(.a(buffered_input), .b(12'b010000010011), .eq(weq1043));
    equaln #(12) e1044(.a(buffered_input), .b(12'b010000010100), .eq(weq1044));
    equaln #(12) e1045(.a(buffered_input), .b(12'b010000010101), .eq(weq1045));
    equaln #(12) e1046(.a(buffered_input), .b(12'b010000010110), .eq(weq1046));
    equaln #(12) e1047(.a(buffered_input), .b(12'b010000010111), .eq(weq1047));
    equaln #(12) e1048(.a(buffered_input), .b(12'b010000011000), .eq(weq1048));
    equaln #(12) e1049(.a(buffered_input), .b(12'b010000011001), .eq(weq1049));
    equaln #(12) e1050(.a(buffered_input), .b(12'b010000011010), .eq(weq1050));
    equaln #(12) e1051(.a(buffered_input), .b(12'b010000011011), .eq(weq1051));
    equaln #(12) e1052(.a(buffered_input), .b(12'b010000011100), .eq(weq1052));
    equaln #(12) e1053(.a(buffered_input), .b(12'b010000011101), .eq(weq1053));
    equaln #(12) e1054(.a(buffered_input), .b(12'b010000011110), .eq(weq1054));
    equaln #(12) e1055(.a(buffered_input), .b(12'b010000011111), .eq(weq1055));
    equaln #(12) e1056(.a(buffered_input), .b(12'b010000100000), .eq(weq1056));
    equaln #(12) e1057(.a(buffered_input), .b(12'b010000100001), .eq(weq1057));
    equaln #(12) e1058(.a(buffered_input), .b(12'b010000100010), .eq(weq1058));
    equaln #(12) e1059(.a(buffered_input), .b(12'b010000100011), .eq(weq1059));
    equaln #(12) e1060(.a(buffered_input), .b(12'b010000100100), .eq(weq1060));
    equaln #(12) e1061(.a(buffered_input), .b(12'b010000100101), .eq(weq1061));
    equaln #(12) e1062(.a(buffered_input), .b(12'b010000100110), .eq(weq1062));
    equaln #(12) e1063(.a(buffered_input), .b(12'b010000100111), .eq(weq1063));
    equaln #(12) e1064(.a(buffered_input), .b(12'b010000101000), .eq(weq1064));
    equaln #(12) e1065(.a(buffered_input), .b(12'b010000101001), .eq(weq1065));
    equaln #(12) e1066(.a(buffered_input), .b(12'b010000101010), .eq(weq1066));
    equaln #(12) e1067(.a(buffered_input), .b(12'b010000101011), .eq(weq1067));
    equaln #(12) e1068(.a(buffered_input), .b(12'b010000101100), .eq(weq1068));
    equaln #(12) e1069(.a(buffered_input), .b(12'b010000101101), .eq(weq1069));
    equaln #(12) e1070(.a(buffered_input), .b(12'b010000101110), .eq(weq1070));
    equaln #(12) e1071(.a(buffered_input), .b(12'b010000101111), .eq(weq1071));
    equaln #(12) e1072(.a(buffered_input), .b(12'b010000110000), .eq(weq1072));
    equaln #(12) e1073(.a(buffered_input), .b(12'b010000110001), .eq(weq1073));
    equaln #(12) e1074(.a(buffered_input), .b(12'b010000110010), .eq(weq1074));
    equaln #(12) e1075(.a(buffered_input), .b(12'b010000110011), .eq(weq1075));
    equaln #(12) e1076(.a(buffered_input), .b(12'b010000110100), .eq(weq1076));
    equaln #(12) e1077(.a(buffered_input), .b(12'b010000110101), .eq(weq1077));
    equaln #(12) e1078(.a(buffered_input), .b(12'b010000110110), .eq(weq1078));
    equaln #(12) e1079(.a(buffered_input), .b(12'b010000110111), .eq(weq1079));
    equaln #(12) e1080(.a(buffered_input), .b(12'b010000111000), .eq(weq1080));
    equaln #(12) e1081(.a(buffered_input), .b(12'b010000111001), .eq(weq1081));
    equaln #(12) e1082(.a(buffered_input), .b(12'b010000111010), .eq(weq1082));
    equaln #(12) e1083(.a(buffered_input), .b(12'b010000111011), .eq(weq1083));
    equaln #(12) e1084(.a(buffered_input), .b(12'b010000111100), .eq(weq1084));
    equaln #(12) e1085(.a(buffered_input), .b(12'b010000111101), .eq(weq1085));
    equaln #(12) e1086(.a(buffered_input), .b(12'b010000111110), .eq(weq1086));
    equaln #(12) e1087(.a(buffered_input), .b(12'b010000111111), .eq(weq1087));
    equaln #(12) e1088(.a(buffered_input), .b(12'b010001000000), .eq(weq1088));
    equaln #(12) e1089(.a(buffered_input), .b(12'b010001000001), .eq(weq1089));
    equaln #(12) e1090(.a(buffered_input), .b(12'b010001000010), .eq(weq1090));
    equaln #(12) e1091(.a(buffered_input), .b(12'b010001000011), .eq(weq1091));
    equaln #(12) e1092(.a(buffered_input), .b(12'b010001000100), .eq(weq1092));
    equaln #(12) e1093(.a(buffered_input), .b(12'b010001000101), .eq(weq1093));
    equaln #(12) e1094(.a(buffered_input), .b(12'b010001000110), .eq(weq1094));
    equaln #(12) e1095(.a(buffered_input), .b(12'b010001000111), .eq(weq1095));
    equaln #(12) e1096(.a(buffered_input), .b(12'b010001001000), .eq(weq1096));
    equaln #(12) e1097(.a(buffered_input), .b(12'b010001001001), .eq(weq1097));
    equaln #(12) e1098(.a(buffered_input), .b(12'b010001001010), .eq(weq1098));
    equaln #(12) e1099(.a(buffered_input), .b(12'b010001001011), .eq(weq1099));
    equaln #(12) e1100(.a(buffered_input), .b(12'b010001001100), .eq(weq1100));
    equaln #(12) e1101(.a(buffered_input), .b(12'b010001001101), .eq(weq1101));
    equaln #(12) e1102(.a(buffered_input), .b(12'b010001001110), .eq(weq1102));
    equaln #(12) e1103(.a(buffered_input), .b(12'b010001001111), .eq(weq1103));
    equaln #(12) e1104(.a(buffered_input), .b(12'b010001010000), .eq(weq1104));
    equaln #(12) e1105(.a(buffered_input), .b(12'b010001010001), .eq(weq1105));
    equaln #(12) e1106(.a(buffered_input), .b(12'b010001010010), .eq(weq1106));
    equaln #(12) e1107(.a(buffered_input), .b(12'b010001010011), .eq(weq1107));
    equaln #(12) e1108(.a(buffered_input), .b(12'b010001010100), .eq(weq1108));
    equaln #(12) e1109(.a(buffered_input), .b(12'b010001010101), .eq(weq1109));
    equaln #(12) e1110(.a(buffered_input), .b(12'b010001010110), .eq(weq1110));
    equaln #(12) e1111(.a(buffered_input), .b(12'b010001010111), .eq(weq1111));
    equaln #(12) e1112(.a(buffered_input), .b(12'b010001011000), .eq(weq1112));
    equaln #(12) e1113(.a(buffered_input), .b(12'b010001011001), .eq(weq1113));
    equaln #(12) e1114(.a(buffered_input), .b(12'b010001011010), .eq(weq1114));
    equaln #(12) e1115(.a(buffered_input), .b(12'b010001011011), .eq(weq1115));
    equaln #(12) e1116(.a(buffered_input), .b(12'b010001011100), .eq(weq1116));
    equaln #(12) e1117(.a(buffered_input), .b(12'b010001011101), .eq(weq1117));
    equaln #(12) e1118(.a(buffered_input), .b(12'b010001011110), .eq(weq1118));
    equaln #(12) e1119(.a(buffered_input), .b(12'b010001011111), .eq(weq1119));
    equaln #(12) e1120(.a(buffered_input), .b(12'b010001100000), .eq(weq1120));
    equaln #(12) e1121(.a(buffered_input), .b(12'b010001100001), .eq(weq1121));
    equaln #(12) e1122(.a(buffered_input), .b(12'b010001100010), .eq(weq1122));
    equaln #(12) e1123(.a(buffered_input), .b(12'b010001100011), .eq(weq1123));
    equaln #(12) e1124(.a(buffered_input), .b(12'b010001100100), .eq(weq1124));
    equaln #(12) e1125(.a(buffered_input), .b(12'b010001100101), .eq(weq1125));
    equaln #(12) e1126(.a(buffered_input), .b(12'b010001100110), .eq(weq1126));
    equaln #(12) e1127(.a(buffered_input), .b(12'b010001100111), .eq(weq1127));
    equaln #(12) e1128(.a(buffered_input), .b(12'b010001101000), .eq(weq1128));
    equaln #(12) e1129(.a(buffered_input), .b(12'b010001101001), .eq(weq1129));
    equaln #(12) e1130(.a(buffered_input), .b(12'b010001101010), .eq(weq1130));
    equaln #(12) e1131(.a(buffered_input), .b(12'b010001101011), .eq(weq1131));
    equaln #(12) e1132(.a(buffered_input), .b(12'b010001101100), .eq(weq1132));
    equaln #(12) e1133(.a(buffered_input), .b(12'b010001101101), .eq(weq1133));
    equaln #(12) e1134(.a(buffered_input), .b(12'b010001101110), .eq(weq1134));
    equaln #(12) e1135(.a(buffered_input), .b(12'b010001101111), .eq(weq1135));
    equaln #(12) e1136(.a(buffered_input), .b(12'b010001110000), .eq(weq1136));
    equaln #(12) e1137(.a(buffered_input), .b(12'b010001110001), .eq(weq1137));
    equaln #(12) e1138(.a(buffered_input), .b(12'b010001110010), .eq(weq1138));
    equaln #(12) e1139(.a(buffered_input), .b(12'b010001110011), .eq(weq1139));
    equaln #(12) e1140(.a(buffered_input), .b(12'b010001110100), .eq(weq1140));
    equaln #(12) e1141(.a(buffered_input), .b(12'b010001110101), .eq(weq1141));
    equaln #(12) e1142(.a(buffered_input), .b(12'b010001110110), .eq(weq1142));
    equaln #(12) e1143(.a(buffered_input), .b(12'b010001110111), .eq(weq1143));
    equaln #(12) e1144(.a(buffered_input), .b(12'b010001111000), .eq(weq1144));
    equaln #(12) e1145(.a(buffered_input), .b(12'b010001111001), .eq(weq1145));
    equaln #(12) e1146(.a(buffered_input), .b(12'b010001111010), .eq(weq1146));
    equaln #(12) e1147(.a(buffered_input), .b(12'b010001111011), .eq(weq1147));
    equaln #(12) e1148(.a(buffered_input), .b(12'b010001111100), .eq(weq1148));
    equaln #(12) e1149(.a(buffered_input), .b(12'b010001111101), .eq(weq1149));
    equaln #(12) e1150(.a(buffered_input), .b(12'b010001111110), .eq(weq1150));
    equaln #(12) e1151(.a(buffered_input), .b(12'b010001111111), .eq(weq1151));
    equaln #(12) e1152(.a(buffered_input), .b(12'b010010000000), .eq(weq1152));
    equaln #(12) e1153(.a(buffered_input), .b(12'b010010000001), .eq(weq1153));
    equaln #(12) e1154(.a(buffered_input), .b(12'b010010000010), .eq(weq1154));
    equaln #(12) e1155(.a(buffered_input), .b(12'b010010000011), .eq(weq1155));
    equaln #(12) e1156(.a(buffered_input), .b(12'b010010000100), .eq(weq1156));
    equaln #(12) e1157(.a(buffered_input), .b(12'b010010000101), .eq(weq1157));
    equaln #(12) e1158(.a(buffered_input), .b(12'b010010000110), .eq(weq1158));
    equaln #(12) e1159(.a(buffered_input), .b(12'b010010000111), .eq(weq1159));
    equaln #(12) e1160(.a(buffered_input), .b(12'b010010001000), .eq(weq1160));
    equaln #(12) e1161(.a(buffered_input), .b(12'b010010001001), .eq(weq1161));
    equaln #(12) e1162(.a(buffered_input), .b(12'b010010001010), .eq(weq1162));
    equaln #(12) e1163(.a(buffered_input), .b(12'b010010001011), .eq(weq1163));
    equaln #(12) e1164(.a(buffered_input), .b(12'b010010001100), .eq(weq1164));
    equaln #(12) e1165(.a(buffered_input), .b(12'b010010001101), .eq(weq1165));
    equaln #(12) e1166(.a(buffered_input), .b(12'b010010001110), .eq(weq1166));
    equaln #(12) e1167(.a(buffered_input), .b(12'b010010001111), .eq(weq1167));
    equaln #(12) e1168(.a(buffered_input), .b(12'b010010010000), .eq(weq1168));
    equaln #(12) e1169(.a(buffered_input), .b(12'b010010010001), .eq(weq1169));
    equaln #(12) e1170(.a(buffered_input), .b(12'b010010010010), .eq(weq1170));
    equaln #(12) e1171(.a(buffered_input), .b(12'b010010010011), .eq(weq1171));
    equaln #(12) e1172(.a(buffered_input), .b(12'b010010010100), .eq(weq1172));
    equaln #(12) e1173(.a(buffered_input), .b(12'b010010010101), .eq(weq1173));
    equaln #(12) e1174(.a(buffered_input), .b(12'b010010010110), .eq(weq1174));
    equaln #(12) e1175(.a(buffered_input), .b(12'b010010010111), .eq(weq1175));
    equaln #(12) e1176(.a(buffered_input), .b(12'b010010011000), .eq(weq1176));
    equaln #(12) e1177(.a(buffered_input), .b(12'b010010011001), .eq(weq1177));
    equaln #(12) e1178(.a(buffered_input), .b(12'b010010011010), .eq(weq1178));
    equaln #(12) e1179(.a(buffered_input), .b(12'b010010011011), .eq(weq1179));
    equaln #(12) e1180(.a(buffered_input), .b(12'b010010011100), .eq(weq1180));
    equaln #(12) e1181(.a(buffered_input), .b(12'b010010011101), .eq(weq1181));
    equaln #(12) e1182(.a(buffered_input), .b(12'b010010011110), .eq(weq1182));
    equaln #(12) e1183(.a(buffered_input), .b(12'b010010011111), .eq(weq1183));
    equaln #(12) e1184(.a(buffered_input), .b(12'b010010100000), .eq(weq1184));
    equaln #(12) e1185(.a(buffered_input), .b(12'b010010100001), .eq(weq1185));
    equaln #(12) e1186(.a(buffered_input), .b(12'b010010100010), .eq(weq1186));
    equaln #(12) e1187(.a(buffered_input), .b(12'b010010100011), .eq(weq1187));
    equaln #(12) e1188(.a(buffered_input), .b(12'b010010100100), .eq(weq1188));
    equaln #(12) e1189(.a(buffered_input), .b(12'b010010100101), .eq(weq1189));
    equaln #(12) e1190(.a(buffered_input), .b(12'b010010100110), .eq(weq1190));
    equaln #(12) e1191(.a(buffered_input), .b(12'b010010100111), .eq(weq1191));
    equaln #(12) e1192(.a(buffered_input), .b(12'b010010101000), .eq(weq1192));
    equaln #(12) e1193(.a(buffered_input), .b(12'b010010101001), .eq(weq1193));
    equaln #(12) e1194(.a(buffered_input), .b(12'b010010101010), .eq(weq1194));
    equaln #(12) e1195(.a(buffered_input), .b(12'b010010101011), .eq(weq1195));
    equaln #(12) e1196(.a(buffered_input), .b(12'b010010101100), .eq(weq1196));
    equaln #(12) e1197(.a(buffered_input), .b(12'b010010101101), .eq(weq1197));
    equaln #(12) e1198(.a(buffered_input), .b(12'b010010101110), .eq(weq1198));
    equaln #(12) e1199(.a(buffered_input), .b(12'b010010101111), .eq(weq1199));
    equaln #(12) e1200(.a(buffered_input), .b(12'b010010110000), .eq(weq1200));
    equaln #(12) e1201(.a(buffered_input), .b(12'b010010110001), .eq(weq1201));
    equaln #(12) e1202(.a(buffered_input), .b(12'b010010110010), .eq(weq1202));
    equaln #(12) e1203(.a(buffered_input), .b(12'b010010110011), .eq(weq1203));
    equaln #(12) e1204(.a(buffered_input), .b(12'b010010110100), .eq(weq1204));
    equaln #(12) e1205(.a(buffered_input), .b(12'b010010110101), .eq(weq1205));
    equaln #(12) e1206(.a(buffered_input), .b(12'b010010110110), .eq(weq1206));
    equaln #(12) e1207(.a(buffered_input), .b(12'b010010110111), .eq(weq1207));
    equaln #(12) e1208(.a(buffered_input), .b(12'b010010111000), .eq(weq1208));
    equaln #(12) e1209(.a(buffered_input), .b(12'b010010111001), .eq(weq1209));
    equaln #(12) e1210(.a(buffered_input), .b(12'b010010111010), .eq(weq1210));
    equaln #(12) e1211(.a(buffered_input), .b(12'b010010111011), .eq(weq1211));
    equaln #(12) e1212(.a(buffered_input), .b(12'b010010111100), .eq(weq1212));
    equaln #(12) e1213(.a(buffered_input), .b(12'b010010111101), .eq(weq1213));
    equaln #(12) e1214(.a(buffered_input), .b(12'b010010111110), .eq(weq1214));
    equaln #(12) e1215(.a(buffered_input), .b(12'b010010111111), .eq(weq1215));
    equaln #(12) e1216(.a(buffered_input), .b(12'b010011000000), .eq(weq1216));
    equaln #(12) e1217(.a(buffered_input), .b(12'b010011000001), .eq(weq1217));
    equaln #(12) e1218(.a(buffered_input), .b(12'b010011000010), .eq(weq1218));
    equaln #(12) e1219(.a(buffered_input), .b(12'b010011000011), .eq(weq1219));
    equaln #(12) e1220(.a(buffered_input), .b(12'b010011000100), .eq(weq1220));
    equaln #(12) e1221(.a(buffered_input), .b(12'b010011000101), .eq(weq1221));
    equaln #(12) e1222(.a(buffered_input), .b(12'b010011000110), .eq(weq1222));
    equaln #(12) e1223(.a(buffered_input), .b(12'b010011000111), .eq(weq1223));
    equaln #(12) e1224(.a(buffered_input), .b(12'b010011001000), .eq(weq1224));
    equaln #(12) e1225(.a(buffered_input), .b(12'b010011001001), .eq(weq1225));
    equaln #(12) e1226(.a(buffered_input), .b(12'b010011001010), .eq(weq1226));
    equaln #(12) e1227(.a(buffered_input), .b(12'b010011001011), .eq(weq1227));
    equaln #(12) e1228(.a(buffered_input), .b(12'b010011001100), .eq(weq1228));
    equaln #(12) e1229(.a(buffered_input), .b(12'b010011001101), .eq(weq1229));
    equaln #(12) e1230(.a(buffered_input), .b(12'b010011001110), .eq(weq1230));
    equaln #(12) e1231(.a(buffered_input), .b(12'b010011001111), .eq(weq1231));
    equaln #(12) e1232(.a(buffered_input), .b(12'b010011010000), .eq(weq1232));
    equaln #(12) e1233(.a(buffered_input), .b(12'b010011010001), .eq(weq1233));
    equaln #(12) e1234(.a(buffered_input), .b(12'b010011010010), .eq(weq1234));
    equaln #(12) e1235(.a(buffered_input), .b(12'b010011010011), .eq(weq1235));
    equaln #(12) e1236(.a(buffered_input), .b(12'b010011010100), .eq(weq1236));
    equaln #(12) e1237(.a(buffered_input), .b(12'b010011010101), .eq(weq1237));
    equaln #(12) e1238(.a(buffered_input), .b(12'b010011010110), .eq(weq1238));
    equaln #(12) e1239(.a(buffered_input), .b(12'b010011010111), .eq(weq1239));
    equaln #(12) e1240(.a(buffered_input), .b(12'b010011011000), .eq(weq1240));
    equaln #(12) e1241(.a(buffered_input), .b(12'b010011011001), .eq(weq1241));
    equaln #(12) e1242(.a(buffered_input), .b(12'b010011011010), .eq(weq1242));
    equaln #(12) e1243(.a(buffered_input), .b(12'b010011011011), .eq(weq1243));
    equaln #(12) e1244(.a(buffered_input), .b(12'b010011011100), .eq(weq1244));
    equaln #(12) e1245(.a(buffered_input), .b(12'b010011011101), .eq(weq1245));
    equaln #(12) e1246(.a(buffered_input), .b(12'b010011011110), .eq(weq1246));
    equaln #(12) e1247(.a(buffered_input), .b(12'b010011011111), .eq(weq1247));
    equaln #(12) e1248(.a(buffered_input), .b(12'b010011100000), .eq(weq1248));
    equaln #(12) e1249(.a(buffered_input), .b(12'b010011100001), .eq(weq1249));
    equaln #(12) e1250(.a(buffered_input), .b(12'b010011100010), .eq(weq1250));
    equaln #(12) e1251(.a(buffered_input), .b(12'b010011100011), .eq(weq1251));
    equaln #(12) e1252(.a(buffered_input), .b(12'b010011100100), .eq(weq1252));
    equaln #(12) e1253(.a(buffered_input), .b(12'b010011100101), .eq(weq1253));
    equaln #(12) e1254(.a(buffered_input), .b(12'b010011100110), .eq(weq1254));
    equaln #(12) e1255(.a(buffered_input), .b(12'b010011100111), .eq(weq1255));
    equaln #(12) e1256(.a(buffered_input), .b(12'b010011101000), .eq(weq1256));
    equaln #(12) e1257(.a(buffered_input), .b(12'b010011101001), .eq(weq1257));
    equaln #(12) e1258(.a(buffered_input), .b(12'b010011101010), .eq(weq1258));
    equaln #(12) e1259(.a(buffered_input), .b(12'b010011101011), .eq(weq1259));
    equaln #(12) e1260(.a(buffered_input), .b(12'b010011101100), .eq(weq1260));
    equaln #(12) e1261(.a(buffered_input), .b(12'b010011101101), .eq(weq1261));
    equaln #(12) e1262(.a(buffered_input), .b(12'b010011101110), .eq(weq1262));
    equaln #(12) e1263(.a(buffered_input), .b(12'b010011101111), .eq(weq1263));
    equaln #(12) e1264(.a(buffered_input), .b(12'b010011110000), .eq(weq1264));
    equaln #(12) e1265(.a(buffered_input), .b(12'b010011110001), .eq(weq1265));
    equaln #(12) e1266(.a(buffered_input), .b(12'b010011110010), .eq(weq1266));
    equaln #(12) e1267(.a(buffered_input), .b(12'b010011110011), .eq(weq1267));
    equaln #(12) e1268(.a(buffered_input), .b(12'b010011110100), .eq(weq1268));
    equaln #(12) e1269(.a(buffered_input), .b(12'b010011110101), .eq(weq1269));
    equaln #(12) e1270(.a(buffered_input), .b(12'b010011110110), .eq(weq1270));
    equaln #(12) e1271(.a(buffered_input), .b(12'b010011110111), .eq(weq1271));
    equaln #(12) e1272(.a(buffered_input), .b(12'b010011111000), .eq(weq1272));
    equaln #(12) e1273(.a(buffered_input), .b(12'b010011111001), .eq(weq1273));
    equaln #(12) e1274(.a(buffered_input), .b(12'b010011111010), .eq(weq1274));
    equaln #(12) e1275(.a(buffered_input), .b(12'b010011111011), .eq(weq1275));
    equaln #(12) e1276(.a(buffered_input), .b(12'b010011111100), .eq(weq1276));
    equaln #(12) e1277(.a(buffered_input), .b(12'b010011111101), .eq(weq1277));
    equaln #(12) e1278(.a(buffered_input), .b(12'b010011111110), .eq(weq1278));
    equaln #(12) e1279(.a(buffered_input), .b(12'b010011111111), .eq(weq1279));
    equaln #(12) e1280(.a(buffered_input), .b(12'b010100000000), .eq(weq1280));
    equaln #(12) e1281(.a(buffered_input), .b(12'b010100000001), .eq(weq1281));
    equaln #(12) e1282(.a(buffered_input), .b(12'b010100000010), .eq(weq1282));
    equaln #(12) e1283(.a(buffered_input), .b(12'b010100000011), .eq(weq1283));
    equaln #(12) e1284(.a(buffered_input), .b(12'b010100000100), .eq(weq1284));
    equaln #(12) e1285(.a(buffered_input), .b(12'b010100000101), .eq(weq1285));
    equaln #(12) e1286(.a(buffered_input), .b(12'b010100000110), .eq(weq1286));
    equaln #(12) e1287(.a(buffered_input), .b(12'b010100000111), .eq(weq1287));
    equaln #(12) e1288(.a(buffered_input), .b(12'b010100001000), .eq(weq1288));
    equaln #(12) e1289(.a(buffered_input), .b(12'b010100001001), .eq(weq1289));
    equaln #(12) e1290(.a(buffered_input), .b(12'b010100001010), .eq(weq1290));
    equaln #(12) e1291(.a(buffered_input), .b(12'b010100001011), .eq(weq1291));
    equaln #(12) e1292(.a(buffered_input), .b(12'b010100001100), .eq(weq1292));
    equaln #(12) e1293(.a(buffered_input), .b(12'b010100001101), .eq(weq1293));
    equaln #(12) e1294(.a(buffered_input), .b(12'b010100001110), .eq(weq1294));
    equaln #(12) e1295(.a(buffered_input), .b(12'b010100001111), .eq(weq1295));
    equaln #(12) e1296(.a(buffered_input), .b(12'b010100010000), .eq(weq1296));
    equaln #(12) e1297(.a(buffered_input), .b(12'b010100010001), .eq(weq1297));
    equaln #(12) e1298(.a(buffered_input), .b(12'b010100010010), .eq(weq1298));
    equaln #(12) e1299(.a(buffered_input), .b(12'b010100010011), .eq(weq1299));
    equaln #(12) e1300(.a(buffered_input), .b(12'b010100010100), .eq(weq1300));
    equaln #(12) e1301(.a(buffered_input), .b(12'b010100010101), .eq(weq1301));
    equaln #(12) e1302(.a(buffered_input), .b(12'b010100010110), .eq(weq1302));
    equaln #(12) e1303(.a(buffered_input), .b(12'b010100010111), .eq(weq1303));
    equaln #(12) e1304(.a(buffered_input), .b(12'b010100011000), .eq(weq1304));
    equaln #(12) e1305(.a(buffered_input), .b(12'b010100011001), .eq(weq1305));
    equaln #(12) e1306(.a(buffered_input), .b(12'b010100011010), .eq(weq1306));
    equaln #(12) e1307(.a(buffered_input), .b(12'b010100011011), .eq(weq1307));
    equaln #(12) e1308(.a(buffered_input), .b(12'b010100011100), .eq(weq1308));
    equaln #(12) e1309(.a(buffered_input), .b(12'b010100011101), .eq(weq1309));
    equaln #(12) e1310(.a(buffered_input), .b(12'b010100011110), .eq(weq1310));
    equaln #(12) e1311(.a(buffered_input), .b(12'b010100011111), .eq(weq1311));
    equaln #(12) e1312(.a(buffered_input), .b(12'b010100100000), .eq(weq1312));
    equaln #(12) e1313(.a(buffered_input), .b(12'b010100100001), .eq(weq1313));
    equaln #(12) e1314(.a(buffered_input), .b(12'b010100100010), .eq(weq1314));
    equaln #(12) e1315(.a(buffered_input), .b(12'b010100100011), .eq(weq1315));
    equaln #(12) e1316(.a(buffered_input), .b(12'b010100100100), .eq(weq1316));
    equaln #(12) e1317(.a(buffered_input), .b(12'b010100100101), .eq(weq1317));
    equaln #(12) e1318(.a(buffered_input), .b(12'b010100100110), .eq(weq1318));
    equaln #(12) e1319(.a(buffered_input), .b(12'b010100100111), .eq(weq1319));
    equaln #(12) e1320(.a(buffered_input), .b(12'b010100101000), .eq(weq1320));
    equaln #(12) e1321(.a(buffered_input), .b(12'b010100101001), .eq(weq1321));
    equaln #(12) e1322(.a(buffered_input), .b(12'b010100101010), .eq(weq1322));
    equaln #(12) e1323(.a(buffered_input), .b(12'b010100101011), .eq(weq1323));
    equaln #(12) e1324(.a(buffered_input), .b(12'b010100101100), .eq(weq1324));
    equaln #(12) e1325(.a(buffered_input), .b(12'b010100101101), .eq(weq1325));
    equaln #(12) e1326(.a(buffered_input), .b(12'b010100101110), .eq(weq1326));
    equaln #(12) e1327(.a(buffered_input), .b(12'b010100101111), .eq(weq1327));
    equaln #(12) e1328(.a(buffered_input), .b(12'b010100110000), .eq(weq1328));
    equaln #(12) e1329(.a(buffered_input), .b(12'b010100110001), .eq(weq1329));
    equaln #(12) e1330(.a(buffered_input), .b(12'b010100110010), .eq(weq1330));
    equaln #(12) e1331(.a(buffered_input), .b(12'b010100110011), .eq(weq1331));
    equaln #(12) e1332(.a(buffered_input), .b(12'b010100110100), .eq(weq1332));
    equaln #(12) e1333(.a(buffered_input), .b(12'b010100110101), .eq(weq1333));
    equaln #(12) e1334(.a(buffered_input), .b(12'b010100110110), .eq(weq1334));
    equaln #(12) e1335(.a(buffered_input), .b(12'b010100110111), .eq(weq1335));
    equaln #(12) e1336(.a(buffered_input), .b(12'b010100111000), .eq(weq1336));
    equaln #(12) e1337(.a(buffered_input), .b(12'b010100111001), .eq(weq1337));
    equaln #(12) e1338(.a(buffered_input), .b(12'b010100111010), .eq(weq1338));
    equaln #(12) e1339(.a(buffered_input), .b(12'b010100111011), .eq(weq1339));
    equaln #(12) e1340(.a(buffered_input), .b(12'b010100111100), .eq(weq1340));
    equaln #(12) e1341(.a(buffered_input), .b(12'b010100111101), .eq(weq1341));
    equaln #(12) e1342(.a(buffered_input), .b(12'b010100111110), .eq(weq1342));
    equaln #(12) e1343(.a(buffered_input), .b(12'b010100111111), .eq(weq1343));
    equaln #(12) e1344(.a(buffered_input), .b(12'b010101000000), .eq(weq1344));
    equaln #(12) e1345(.a(buffered_input), .b(12'b010101000001), .eq(weq1345));
    equaln #(12) e1346(.a(buffered_input), .b(12'b010101000010), .eq(weq1346));
    equaln #(12) e1347(.a(buffered_input), .b(12'b010101000011), .eq(weq1347));
    equaln #(12) e1348(.a(buffered_input), .b(12'b010101000100), .eq(weq1348));
    equaln #(12) e1349(.a(buffered_input), .b(12'b010101000101), .eq(weq1349));
    equaln #(12) e1350(.a(buffered_input), .b(12'b010101000110), .eq(weq1350));
    equaln #(12) e1351(.a(buffered_input), .b(12'b010101000111), .eq(weq1351));
    equaln #(12) e1352(.a(buffered_input), .b(12'b010101001000), .eq(weq1352));
    equaln #(12) e1353(.a(buffered_input), .b(12'b010101001001), .eq(weq1353));
    equaln #(12) e1354(.a(buffered_input), .b(12'b010101001010), .eq(weq1354));
    equaln #(12) e1355(.a(buffered_input), .b(12'b010101001011), .eq(weq1355));
    equaln #(12) e1356(.a(buffered_input), .b(12'b010101001100), .eq(weq1356));
    equaln #(12) e1357(.a(buffered_input), .b(12'b010101001101), .eq(weq1357));
    equaln #(12) e1358(.a(buffered_input), .b(12'b010101001110), .eq(weq1358));
    equaln #(12) e1359(.a(buffered_input), .b(12'b010101001111), .eq(weq1359));
    equaln #(12) e1360(.a(buffered_input), .b(12'b010101010000), .eq(weq1360));
    equaln #(12) e1361(.a(buffered_input), .b(12'b010101010001), .eq(weq1361));
    equaln #(12) e1362(.a(buffered_input), .b(12'b010101010010), .eq(weq1362));
    equaln #(12) e1363(.a(buffered_input), .b(12'b010101010011), .eq(weq1363));
    equaln #(12) e1364(.a(buffered_input), .b(12'b010101010100), .eq(weq1364));
    equaln #(12) e1365(.a(buffered_input), .b(12'b010101010101), .eq(weq1365));
    equaln #(12) e1366(.a(buffered_input), .b(12'b010101010110), .eq(weq1366));
    equaln #(12) e1367(.a(buffered_input), .b(12'b010101010111), .eq(weq1367));
    equaln #(12) e1368(.a(buffered_input), .b(12'b010101011000), .eq(weq1368));
    equaln #(12) e1369(.a(buffered_input), .b(12'b010101011001), .eq(weq1369));
    equaln #(12) e1370(.a(buffered_input), .b(12'b010101011010), .eq(weq1370));
    equaln #(12) e1371(.a(buffered_input), .b(12'b010101011011), .eq(weq1371));
    equaln #(12) e1372(.a(buffered_input), .b(12'b010101011100), .eq(weq1372));
    equaln #(12) e1373(.a(buffered_input), .b(12'b010101011101), .eq(weq1373));
    equaln #(12) e1374(.a(buffered_input), .b(12'b010101011110), .eq(weq1374));
    equaln #(12) e1375(.a(buffered_input), .b(12'b010101011111), .eq(weq1375));
    equaln #(12) e1376(.a(buffered_input), .b(12'b010101100000), .eq(weq1376));
    equaln #(12) e1377(.a(buffered_input), .b(12'b010101100001), .eq(weq1377));
    equaln #(12) e1378(.a(buffered_input), .b(12'b010101100010), .eq(weq1378));
    equaln #(12) e1379(.a(buffered_input), .b(12'b010101100011), .eq(weq1379));
    equaln #(12) e1380(.a(buffered_input), .b(12'b010101100100), .eq(weq1380));
    equaln #(12) e1381(.a(buffered_input), .b(12'b010101100101), .eq(weq1381));
    equaln #(12) e1382(.a(buffered_input), .b(12'b010101100110), .eq(weq1382));
    equaln #(12) e1383(.a(buffered_input), .b(12'b010101100111), .eq(weq1383));
    equaln #(12) e1384(.a(buffered_input), .b(12'b010101101000), .eq(weq1384));
    equaln #(12) e1385(.a(buffered_input), .b(12'b010101101001), .eq(weq1385));
    equaln #(12) e1386(.a(buffered_input), .b(12'b010101101010), .eq(weq1386));
    equaln #(12) e1387(.a(buffered_input), .b(12'b010101101011), .eq(weq1387));
    equaln #(12) e1388(.a(buffered_input), .b(12'b010101101100), .eq(weq1388));
    equaln #(12) e1389(.a(buffered_input), .b(12'b010101101101), .eq(weq1389));
    equaln #(12) e1390(.a(buffered_input), .b(12'b010101101110), .eq(weq1390));
    equaln #(12) e1391(.a(buffered_input), .b(12'b010101101111), .eq(weq1391));
    equaln #(12) e1392(.a(buffered_input), .b(12'b010101110000), .eq(weq1392));
    equaln #(12) e1393(.a(buffered_input), .b(12'b010101110001), .eq(weq1393));
    equaln #(12) e1394(.a(buffered_input), .b(12'b010101110010), .eq(weq1394));
    equaln #(12) e1395(.a(buffered_input), .b(12'b010101110011), .eq(weq1395));
    equaln #(12) e1396(.a(buffered_input), .b(12'b010101110100), .eq(weq1396));
    equaln #(12) e1397(.a(buffered_input), .b(12'b010101110101), .eq(weq1397));
    equaln #(12) e1398(.a(buffered_input), .b(12'b010101110110), .eq(weq1398));
    equaln #(12) e1399(.a(buffered_input), .b(12'b010101110111), .eq(weq1399));
    equaln #(12) e1400(.a(buffered_input), .b(12'b010101111000), .eq(weq1400));
    equaln #(12) e1401(.a(buffered_input), .b(12'b010101111001), .eq(weq1401));
    equaln #(12) e1402(.a(buffered_input), .b(12'b010101111010), .eq(weq1402));
    equaln #(12) e1403(.a(buffered_input), .b(12'b010101111011), .eq(weq1403));
    equaln #(12) e1404(.a(buffered_input), .b(12'b010101111100), .eq(weq1404));
    equaln #(12) e1405(.a(buffered_input), .b(12'b010101111101), .eq(weq1405));
    equaln #(12) e1406(.a(buffered_input), .b(12'b010101111110), .eq(weq1406));
    equaln #(12) e1407(.a(buffered_input), .b(12'b010101111111), .eq(weq1407));
    equaln #(12) e1408(.a(buffered_input), .b(12'b010110000000), .eq(weq1408));
    equaln #(12) e1409(.a(buffered_input), .b(12'b010110000001), .eq(weq1409));
    equaln #(12) e1410(.a(buffered_input), .b(12'b010110000010), .eq(weq1410));
    equaln #(12) e1411(.a(buffered_input), .b(12'b010110000011), .eq(weq1411));
    equaln #(12) e1412(.a(buffered_input), .b(12'b010110000100), .eq(weq1412));
    equaln #(12) e1413(.a(buffered_input), .b(12'b010110000101), .eq(weq1413));
    equaln #(12) e1414(.a(buffered_input), .b(12'b010110000110), .eq(weq1414));
    equaln #(12) e1415(.a(buffered_input), .b(12'b010110000111), .eq(weq1415));
    equaln #(12) e1416(.a(buffered_input), .b(12'b010110001000), .eq(weq1416));
    equaln #(12) e1417(.a(buffered_input), .b(12'b010110001001), .eq(weq1417));
    equaln #(12) e1418(.a(buffered_input), .b(12'b010110001010), .eq(weq1418));
    equaln #(12) e1419(.a(buffered_input), .b(12'b010110001011), .eq(weq1419));
    equaln #(12) e1420(.a(buffered_input), .b(12'b010110001100), .eq(weq1420));
    equaln #(12) e1421(.a(buffered_input), .b(12'b010110001101), .eq(weq1421));
    equaln #(12) e1422(.a(buffered_input), .b(12'b010110001110), .eq(weq1422));
    equaln #(12) e1423(.a(buffered_input), .b(12'b010110001111), .eq(weq1423));
    equaln #(12) e1424(.a(buffered_input), .b(12'b010110010000), .eq(weq1424));
    equaln #(12) e1425(.a(buffered_input), .b(12'b010110010001), .eq(weq1425));
    equaln #(12) e1426(.a(buffered_input), .b(12'b010110010010), .eq(weq1426));
    equaln #(12) e1427(.a(buffered_input), .b(12'b010110010011), .eq(weq1427));
    equaln #(12) e1428(.a(buffered_input), .b(12'b010110010100), .eq(weq1428));
    equaln #(12) e1429(.a(buffered_input), .b(12'b010110010101), .eq(weq1429));
    equaln #(12) e1430(.a(buffered_input), .b(12'b010110010110), .eq(weq1430));
    equaln #(12) e1431(.a(buffered_input), .b(12'b010110010111), .eq(weq1431));
    equaln #(12) e1432(.a(buffered_input), .b(12'b010110011000), .eq(weq1432));
    equaln #(12) e1433(.a(buffered_input), .b(12'b010110011001), .eq(weq1433));
    equaln #(12) e1434(.a(buffered_input), .b(12'b010110011010), .eq(weq1434));
    equaln #(12) e1435(.a(buffered_input), .b(12'b010110011011), .eq(weq1435));
    equaln #(12) e1436(.a(buffered_input), .b(12'b010110011100), .eq(weq1436));
    equaln #(12) e1437(.a(buffered_input), .b(12'b010110011101), .eq(weq1437));
    equaln #(12) e1438(.a(buffered_input), .b(12'b010110011110), .eq(weq1438));
    equaln #(12) e1439(.a(buffered_input), .b(12'b010110011111), .eq(weq1439));
    equaln #(12) e1440(.a(buffered_input), .b(12'b010110100000), .eq(weq1440));
    equaln #(12) e1441(.a(buffered_input), .b(12'b010110100001), .eq(weq1441));
    equaln #(12) e1442(.a(buffered_input), .b(12'b010110100010), .eq(weq1442));
    equaln #(12) e1443(.a(buffered_input), .b(12'b010110100011), .eq(weq1443));
    equaln #(12) e1444(.a(buffered_input), .b(12'b010110100100), .eq(weq1444));
    equaln #(12) e1445(.a(buffered_input), .b(12'b010110100101), .eq(weq1445));
    equaln #(12) e1446(.a(buffered_input), .b(12'b010110100110), .eq(weq1446));
    equaln #(12) e1447(.a(buffered_input), .b(12'b010110100111), .eq(weq1447));
    equaln #(12) e1448(.a(buffered_input), .b(12'b010110101000), .eq(weq1448));
    equaln #(12) e1449(.a(buffered_input), .b(12'b010110101001), .eq(weq1449));
    equaln #(12) e1450(.a(buffered_input), .b(12'b010110101010), .eq(weq1450));
    equaln #(12) e1451(.a(buffered_input), .b(12'b010110101011), .eq(weq1451));
    equaln #(12) e1452(.a(buffered_input), .b(12'b010110101100), .eq(weq1452));
    equaln #(12) e1453(.a(buffered_input), .b(12'b010110101101), .eq(weq1453));
    equaln #(12) e1454(.a(buffered_input), .b(12'b010110101110), .eq(weq1454));
    equaln #(12) e1455(.a(buffered_input), .b(12'b010110101111), .eq(weq1455));
    equaln #(12) e1456(.a(buffered_input), .b(12'b010110110000), .eq(weq1456));
    equaln #(12) e1457(.a(buffered_input), .b(12'b010110110001), .eq(weq1457));
    equaln #(12) e1458(.a(buffered_input), .b(12'b010110110010), .eq(weq1458));
    equaln #(12) e1459(.a(buffered_input), .b(12'b010110110011), .eq(weq1459));
    equaln #(12) e1460(.a(buffered_input), .b(12'b010110110100), .eq(weq1460));
    equaln #(12) e1461(.a(buffered_input), .b(12'b010110110101), .eq(weq1461));
    equaln #(12) e1462(.a(buffered_input), .b(12'b010110110110), .eq(weq1462));
    equaln #(12) e1463(.a(buffered_input), .b(12'b010110110111), .eq(weq1463));
    equaln #(12) e1464(.a(buffered_input), .b(12'b010110111000), .eq(weq1464));
    equaln #(12) e1465(.a(buffered_input), .b(12'b010110111001), .eq(weq1465));
    equaln #(12) e1466(.a(buffered_input), .b(12'b010110111010), .eq(weq1466));
    equaln #(12) e1467(.a(buffered_input), .b(12'b010110111011), .eq(weq1467));
    equaln #(12) e1468(.a(buffered_input), .b(12'b010110111100), .eq(weq1468));
    equaln #(12) e1469(.a(buffered_input), .b(12'b010110111101), .eq(weq1469));
    equaln #(12) e1470(.a(buffered_input), .b(12'b010110111110), .eq(weq1470));
    equaln #(12) e1471(.a(buffered_input), .b(12'b010110111111), .eq(weq1471));
    equaln #(12) e1472(.a(buffered_input), .b(12'b010111000000), .eq(weq1472));
    equaln #(12) e1473(.a(buffered_input), .b(12'b010111000001), .eq(weq1473));
    equaln #(12) e1474(.a(buffered_input), .b(12'b010111000010), .eq(weq1474));
    equaln #(12) e1475(.a(buffered_input), .b(12'b010111000011), .eq(weq1475));
    equaln #(12) e1476(.a(buffered_input), .b(12'b010111000100), .eq(weq1476));
    equaln #(12) e1477(.a(buffered_input), .b(12'b010111000101), .eq(weq1477));
    equaln #(12) e1478(.a(buffered_input), .b(12'b010111000110), .eq(weq1478));
    equaln #(12) e1479(.a(buffered_input), .b(12'b010111000111), .eq(weq1479));
    equaln #(12) e1480(.a(buffered_input), .b(12'b010111001000), .eq(weq1480));
    equaln #(12) e1481(.a(buffered_input), .b(12'b010111001001), .eq(weq1481));
    equaln #(12) e1482(.a(buffered_input), .b(12'b010111001010), .eq(weq1482));
    equaln #(12) e1483(.a(buffered_input), .b(12'b010111001011), .eq(weq1483));
    equaln #(12) e1484(.a(buffered_input), .b(12'b010111001100), .eq(weq1484));
    equaln #(12) e1485(.a(buffered_input), .b(12'b010111001101), .eq(weq1485));
    equaln #(12) e1486(.a(buffered_input), .b(12'b010111001110), .eq(weq1486));
    equaln #(12) e1487(.a(buffered_input), .b(12'b010111001111), .eq(weq1487));
    equaln #(12) e1488(.a(buffered_input), .b(12'b010111010000), .eq(weq1488));
    equaln #(12) e1489(.a(buffered_input), .b(12'b010111010001), .eq(weq1489));
    equaln #(12) e1490(.a(buffered_input), .b(12'b010111010010), .eq(weq1490));
    equaln #(12) e1491(.a(buffered_input), .b(12'b010111010011), .eq(weq1491));
    equaln #(12) e1492(.a(buffered_input), .b(12'b010111010100), .eq(weq1492));
    equaln #(12) e1493(.a(buffered_input), .b(12'b010111010101), .eq(weq1493));
    equaln #(12) e1494(.a(buffered_input), .b(12'b010111010110), .eq(weq1494));
    equaln #(12) e1495(.a(buffered_input), .b(12'b010111010111), .eq(weq1495));
    equaln #(12) e1496(.a(buffered_input), .b(12'b010111011000), .eq(weq1496));
    equaln #(12) e1497(.a(buffered_input), .b(12'b010111011001), .eq(weq1497));
    equaln #(12) e1498(.a(buffered_input), .b(12'b010111011010), .eq(weq1498));
    equaln #(12) e1499(.a(buffered_input), .b(12'b010111011011), .eq(weq1499));
    equaln #(12) e1500(.a(buffered_input), .b(12'b010111011100), .eq(weq1500));
    equaln #(12) e1501(.a(buffered_input), .b(12'b010111011101), .eq(weq1501));
    equaln #(12) e1502(.a(buffered_input), .b(12'b010111011110), .eq(weq1502));
    equaln #(12) e1503(.a(buffered_input), .b(12'b010111011111), .eq(weq1503));
    equaln #(12) e1504(.a(buffered_input), .b(12'b010111100000), .eq(weq1504));
    equaln #(12) e1505(.a(buffered_input), .b(12'b010111100001), .eq(weq1505));
    equaln #(12) e1506(.a(buffered_input), .b(12'b010111100010), .eq(weq1506));
    equaln #(12) e1507(.a(buffered_input), .b(12'b010111100011), .eq(weq1507));
    equaln #(12) e1508(.a(buffered_input), .b(12'b010111100100), .eq(weq1508));
    equaln #(12) e1509(.a(buffered_input), .b(12'b010111100101), .eq(weq1509));
    equaln #(12) e1510(.a(buffered_input), .b(12'b010111100110), .eq(weq1510));
    equaln #(12) e1511(.a(buffered_input), .b(12'b010111100111), .eq(weq1511));
    equaln #(12) e1512(.a(buffered_input), .b(12'b010111101000), .eq(weq1512));
    equaln #(12) e1513(.a(buffered_input), .b(12'b010111101001), .eq(weq1513));
    equaln #(12) e1514(.a(buffered_input), .b(12'b010111101010), .eq(weq1514));
    equaln #(12) e1515(.a(buffered_input), .b(12'b010111101011), .eq(weq1515));
    equaln #(12) e1516(.a(buffered_input), .b(12'b010111101100), .eq(weq1516));
    equaln #(12) e1517(.a(buffered_input), .b(12'b010111101101), .eq(weq1517));
    equaln #(12) e1518(.a(buffered_input), .b(12'b010111101110), .eq(weq1518));
    equaln #(12) e1519(.a(buffered_input), .b(12'b010111101111), .eq(weq1519));
    equaln #(12) e1520(.a(buffered_input), .b(12'b010111110000), .eq(weq1520));
    equaln #(12) e1521(.a(buffered_input), .b(12'b010111110001), .eq(weq1521));
    equaln #(12) e1522(.a(buffered_input), .b(12'b010111110010), .eq(weq1522));
    equaln #(12) e1523(.a(buffered_input), .b(12'b010111110011), .eq(weq1523));
    equaln #(12) e1524(.a(buffered_input), .b(12'b010111110100), .eq(weq1524));
    equaln #(12) e1525(.a(buffered_input), .b(12'b010111110101), .eq(weq1525));
    equaln #(12) e1526(.a(buffered_input), .b(12'b010111110110), .eq(weq1526));
    equaln #(12) e1527(.a(buffered_input), .b(12'b010111110111), .eq(weq1527));
    equaln #(12) e1528(.a(buffered_input), .b(12'b010111111000), .eq(weq1528));
    equaln #(12) e1529(.a(buffered_input), .b(12'b010111111001), .eq(weq1529));
    equaln #(12) e1530(.a(buffered_input), .b(12'b010111111010), .eq(weq1530));
    equaln #(12) e1531(.a(buffered_input), .b(12'b010111111011), .eq(weq1531));
    equaln #(12) e1532(.a(buffered_input), .b(12'b010111111100), .eq(weq1532));
    equaln #(12) e1533(.a(buffered_input), .b(12'b010111111101), .eq(weq1533));
    equaln #(12) e1534(.a(buffered_input), .b(12'b010111111110), .eq(weq1534));
    equaln #(12) e1535(.a(buffered_input), .b(12'b010111111111), .eq(weq1535));
    equaln #(12) e1536(.a(buffered_input), .b(12'b011000000000), .eq(weq1536));
    equaln #(12) e1537(.a(buffered_input), .b(12'b011000000001), .eq(weq1537));
    equaln #(12) e1538(.a(buffered_input), .b(12'b011000000010), .eq(weq1538));
    equaln #(12) e1539(.a(buffered_input), .b(12'b011000000011), .eq(weq1539));
    equaln #(12) e1540(.a(buffered_input), .b(12'b011000000100), .eq(weq1540));
    equaln #(12) e1541(.a(buffered_input), .b(12'b011000000101), .eq(weq1541));
    equaln #(12) e1542(.a(buffered_input), .b(12'b011000000110), .eq(weq1542));
    equaln #(12) e1543(.a(buffered_input), .b(12'b011000000111), .eq(weq1543));
    equaln #(12) e1544(.a(buffered_input), .b(12'b011000001000), .eq(weq1544));
    equaln #(12) e1545(.a(buffered_input), .b(12'b011000001001), .eq(weq1545));
    equaln #(12) e1546(.a(buffered_input), .b(12'b011000001010), .eq(weq1546));
    equaln #(12) e1547(.a(buffered_input), .b(12'b011000001011), .eq(weq1547));
    equaln #(12) e1548(.a(buffered_input), .b(12'b011000001100), .eq(weq1548));
    equaln #(12) e1549(.a(buffered_input), .b(12'b011000001101), .eq(weq1549));
    equaln #(12) e1550(.a(buffered_input), .b(12'b011000001110), .eq(weq1550));
    equaln #(12) e1551(.a(buffered_input), .b(12'b011000001111), .eq(weq1551));
    equaln #(12) e1552(.a(buffered_input), .b(12'b011000010000), .eq(weq1552));
    equaln #(12) e1553(.a(buffered_input), .b(12'b011000010001), .eq(weq1553));
    equaln #(12) e1554(.a(buffered_input), .b(12'b011000010010), .eq(weq1554));
    equaln #(12) e1555(.a(buffered_input), .b(12'b011000010011), .eq(weq1555));
    equaln #(12) e1556(.a(buffered_input), .b(12'b011000010100), .eq(weq1556));
    equaln #(12) e1557(.a(buffered_input), .b(12'b011000010101), .eq(weq1557));
    equaln #(12) e1558(.a(buffered_input), .b(12'b011000010110), .eq(weq1558));
    equaln #(12) e1559(.a(buffered_input), .b(12'b011000010111), .eq(weq1559));
    equaln #(12) e1560(.a(buffered_input), .b(12'b011000011000), .eq(weq1560));
    equaln #(12) e1561(.a(buffered_input), .b(12'b011000011001), .eq(weq1561));
    equaln #(12) e1562(.a(buffered_input), .b(12'b011000011010), .eq(weq1562));
    equaln #(12) e1563(.a(buffered_input), .b(12'b011000011011), .eq(weq1563));
    equaln #(12) e1564(.a(buffered_input), .b(12'b011000011100), .eq(weq1564));
    equaln #(12) e1565(.a(buffered_input), .b(12'b011000011101), .eq(weq1565));
    equaln #(12) e1566(.a(buffered_input), .b(12'b011000011110), .eq(weq1566));
    equaln #(12) e1567(.a(buffered_input), .b(12'b011000011111), .eq(weq1567));
    equaln #(12) e1568(.a(buffered_input), .b(12'b011000100000), .eq(weq1568));
    equaln #(12) e1569(.a(buffered_input), .b(12'b011000100001), .eq(weq1569));
    equaln #(12) e1570(.a(buffered_input), .b(12'b011000100010), .eq(weq1570));
    equaln #(12) e1571(.a(buffered_input), .b(12'b011000100011), .eq(weq1571));
    equaln #(12) e1572(.a(buffered_input), .b(12'b011000100100), .eq(weq1572));
    equaln #(12) e1573(.a(buffered_input), .b(12'b011000100101), .eq(weq1573));
    equaln #(12) e1574(.a(buffered_input), .b(12'b011000100110), .eq(weq1574));
    equaln #(12) e1575(.a(buffered_input), .b(12'b011000100111), .eq(weq1575));
    equaln #(12) e1576(.a(buffered_input), .b(12'b011000101000), .eq(weq1576));
    equaln #(12) e1577(.a(buffered_input), .b(12'b011000101001), .eq(weq1577));
    equaln #(12) e1578(.a(buffered_input), .b(12'b011000101010), .eq(weq1578));
    equaln #(12) e1579(.a(buffered_input), .b(12'b011000101011), .eq(weq1579));
    equaln #(12) e1580(.a(buffered_input), .b(12'b011000101100), .eq(weq1580));
    equaln #(12) e1581(.a(buffered_input), .b(12'b011000101101), .eq(weq1581));
    equaln #(12) e1582(.a(buffered_input), .b(12'b011000101110), .eq(weq1582));
    equaln #(12) e1583(.a(buffered_input), .b(12'b011000101111), .eq(weq1583));
    equaln #(12) e1584(.a(buffered_input), .b(12'b011000110000), .eq(weq1584));
    equaln #(12) e1585(.a(buffered_input), .b(12'b011000110001), .eq(weq1585));
    equaln #(12) e1586(.a(buffered_input), .b(12'b011000110010), .eq(weq1586));
    equaln #(12) e1587(.a(buffered_input), .b(12'b011000110011), .eq(weq1587));
    equaln #(12) e1588(.a(buffered_input), .b(12'b011000110100), .eq(weq1588));
    equaln #(12) e1589(.a(buffered_input), .b(12'b011000110101), .eq(weq1589));
    equaln #(12) e1590(.a(buffered_input), .b(12'b011000110110), .eq(weq1590));
    equaln #(12) e1591(.a(buffered_input), .b(12'b011000110111), .eq(weq1591));
    equaln #(12) e1592(.a(buffered_input), .b(12'b011000111000), .eq(weq1592));
    equaln #(12) e1593(.a(buffered_input), .b(12'b011000111001), .eq(weq1593));
    equaln #(12) e1594(.a(buffered_input), .b(12'b011000111010), .eq(weq1594));
    equaln #(12) e1595(.a(buffered_input), .b(12'b011000111011), .eq(weq1595));
    equaln #(12) e1596(.a(buffered_input), .b(12'b011000111100), .eq(weq1596));
    equaln #(12) e1597(.a(buffered_input), .b(12'b011000111101), .eq(weq1597));
    equaln #(12) e1598(.a(buffered_input), .b(12'b011000111110), .eq(weq1598));
    equaln #(12) e1599(.a(buffered_input), .b(12'b011000111111), .eq(weq1599));
    equaln #(12) e1600(.a(buffered_input), .b(12'b011001000000), .eq(weq1600));
    equaln #(12) e1601(.a(buffered_input), .b(12'b011001000001), .eq(weq1601));
    equaln #(12) e1602(.a(buffered_input), .b(12'b011001000010), .eq(weq1602));
    equaln #(12) e1603(.a(buffered_input), .b(12'b011001000011), .eq(weq1603));
    equaln #(12) e1604(.a(buffered_input), .b(12'b011001000100), .eq(weq1604));
    equaln #(12) e1605(.a(buffered_input), .b(12'b011001000101), .eq(weq1605));
    equaln #(12) e1606(.a(buffered_input), .b(12'b011001000110), .eq(weq1606));
    equaln #(12) e1607(.a(buffered_input), .b(12'b011001000111), .eq(weq1607));
    equaln #(12) e1608(.a(buffered_input), .b(12'b011001001000), .eq(weq1608));
    equaln #(12) e1609(.a(buffered_input), .b(12'b011001001001), .eq(weq1609));
    equaln #(12) e1610(.a(buffered_input), .b(12'b011001001010), .eq(weq1610));
    equaln #(12) e1611(.a(buffered_input), .b(12'b011001001011), .eq(weq1611));
    equaln #(12) e1612(.a(buffered_input), .b(12'b011001001100), .eq(weq1612));
    equaln #(12) e1613(.a(buffered_input), .b(12'b011001001101), .eq(weq1613));
    equaln #(12) e1614(.a(buffered_input), .b(12'b011001001110), .eq(weq1614));
    equaln #(12) e1615(.a(buffered_input), .b(12'b011001001111), .eq(weq1615));
    equaln #(12) e1616(.a(buffered_input), .b(12'b011001010000), .eq(weq1616));
    equaln #(12) e1617(.a(buffered_input), .b(12'b011001010001), .eq(weq1617));
    equaln #(12) e1618(.a(buffered_input), .b(12'b011001010010), .eq(weq1618));
    equaln #(12) e1619(.a(buffered_input), .b(12'b011001010011), .eq(weq1619));
    equaln #(12) e1620(.a(buffered_input), .b(12'b011001010100), .eq(weq1620));
    equaln #(12) e1621(.a(buffered_input), .b(12'b011001010101), .eq(weq1621));
    equaln #(12) e1622(.a(buffered_input), .b(12'b011001010110), .eq(weq1622));
    equaln #(12) e1623(.a(buffered_input), .b(12'b011001010111), .eq(weq1623));
    equaln #(12) e1624(.a(buffered_input), .b(12'b011001011000), .eq(weq1624));
    equaln #(12) e1625(.a(buffered_input), .b(12'b011001011001), .eq(weq1625));
    equaln #(12) e1626(.a(buffered_input), .b(12'b011001011010), .eq(weq1626));
    equaln #(12) e1627(.a(buffered_input), .b(12'b011001011011), .eq(weq1627));
    equaln #(12) e1628(.a(buffered_input), .b(12'b011001011100), .eq(weq1628));
    equaln #(12) e1629(.a(buffered_input), .b(12'b011001011101), .eq(weq1629));
    equaln #(12) e1630(.a(buffered_input), .b(12'b011001011110), .eq(weq1630));
    equaln #(12) e1631(.a(buffered_input), .b(12'b011001011111), .eq(weq1631));
    equaln #(12) e1632(.a(buffered_input), .b(12'b011001100000), .eq(weq1632));
    equaln #(12) e1633(.a(buffered_input), .b(12'b011001100001), .eq(weq1633));
    equaln #(12) e1634(.a(buffered_input), .b(12'b011001100010), .eq(weq1634));
    equaln #(12) e1635(.a(buffered_input), .b(12'b011001100011), .eq(weq1635));
    equaln #(12) e1636(.a(buffered_input), .b(12'b011001100100), .eq(weq1636));
    equaln #(12) e1637(.a(buffered_input), .b(12'b011001100101), .eq(weq1637));
    equaln #(12) e1638(.a(buffered_input), .b(12'b011001100110), .eq(weq1638));
    equaln #(12) e1639(.a(buffered_input), .b(12'b011001100111), .eq(weq1639));
    equaln #(12) e1640(.a(buffered_input), .b(12'b011001101000), .eq(weq1640));
    equaln #(12) e1641(.a(buffered_input), .b(12'b011001101001), .eq(weq1641));
    equaln #(12) e1642(.a(buffered_input), .b(12'b011001101010), .eq(weq1642));
    equaln #(12) e1643(.a(buffered_input), .b(12'b011001101011), .eq(weq1643));
    equaln #(12) e1644(.a(buffered_input), .b(12'b011001101100), .eq(weq1644));
    equaln #(12) e1645(.a(buffered_input), .b(12'b011001101101), .eq(weq1645));
    equaln #(12) e1646(.a(buffered_input), .b(12'b011001101110), .eq(weq1646));
    equaln #(12) e1647(.a(buffered_input), .b(12'b011001101111), .eq(weq1647));
    equaln #(12) e1648(.a(buffered_input), .b(12'b011001110000), .eq(weq1648));
    equaln #(12) e1649(.a(buffered_input), .b(12'b011001110001), .eq(weq1649));
    equaln #(12) e1650(.a(buffered_input), .b(12'b011001110010), .eq(weq1650));
    equaln #(12) e1651(.a(buffered_input), .b(12'b011001110011), .eq(weq1651));
    equaln #(12) e1652(.a(buffered_input), .b(12'b011001110100), .eq(weq1652));
    equaln #(12) e1653(.a(buffered_input), .b(12'b011001110101), .eq(weq1653));
    equaln #(12) e1654(.a(buffered_input), .b(12'b011001110110), .eq(weq1654));
    equaln #(12) e1655(.a(buffered_input), .b(12'b011001110111), .eq(weq1655));
    equaln #(12) e1656(.a(buffered_input), .b(12'b011001111000), .eq(weq1656));
    equaln #(12) e1657(.a(buffered_input), .b(12'b011001111001), .eq(weq1657));
    equaln #(12) e1658(.a(buffered_input), .b(12'b011001111010), .eq(weq1658));
    equaln #(12) e1659(.a(buffered_input), .b(12'b011001111011), .eq(weq1659));
    equaln #(12) e1660(.a(buffered_input), .b(12'b011001111100), .eq(weq1660));
    equaln #(12) e1661(.a(buffered_input), .b(12'b011001111101), .eq(weq1661));
    equaln #(12) e1662(.a(buffered_input), .b(12'b011001111110), .eq(weq1662));
    equaln #(12) e1663(.a(buffered_input), .b(12'b011001111111), .eq(weq1663));
    equaln #(12) e1664(.a(buffered_input), .b(12'b011010000000), .eq(weq1664));
    equaln #(12) e1665(.a(buffered_input), .b(12'b011010000001), .eq(weq1665));
    equaln #(12) e1666(.a(buffered_input), .b(12'b011010000010), .eq(weq1666));
    equaln #(12) e1667(.a(buffered_input), .b(12'b011010000011), .eq(weq1667));
    equaln #(12) e1668(.a(buffered_input), .b(12'b011010000100), .eq(weq1668));
    equaln #(12) e1669(.a(buffered_input), .b(12'b011010000101), .eq(weq1669));
    equaln #(12) e1670(.a(buffered_input), .b(12'b011010000110), .eq(weq1670));
    equaln #(12) e1671(.a(buffered_input), .b(12'b011010000111), .eq(weq1671));
    equaln #(12) e1672(.a(buffered_input), .b(12'b011010001000), .eq(weq1672));
    equaln #(12) e1673(.a(buffered_input), .b(12'b011010001001), .eq(weq1673));
    equaln #(12) e1674(.a(buffered_input), .b(12'b011010001010), .eq(weq1674));
    equaln #(12) e1675(.a(buffered_input), .b(12'b011010001011), .eq(weq1675));
    equaln #(12) e1676(.a(buffered_input), .b(12'b011010001100), .eq(weq1676));
    equaln #(12) e1677(.a(buffered_input), .b(12'b011010001101), .eq(weq1677));
    equaln #(12) e1678(.a(buffered_input), .b(12'b011010001110), .eq(weq1678));
    equaln #(12) e1679(.a(buffered_input), .b(12'b011010001111), .eq(weq1679));
    equaln #(12) e1680(.a(buffered_input), .b(12'b011010010000), .eq(weq1680));
    equaln #(12) e1681(.a(buffered_input), .b(12'b011010010001), .eq(weq1681));
    equaln #(12) e1682(.a(buffered_input), .b(12'b011010010010), .eq(weq1682));
    equaln #(12) e1683(.a(buffered_input), .b(12'b011010010011), .eq(weq1683));
    equaln #(12) e1684(.a(buffered_input), .b(12'b011010010100), .eq(weq1684));
    equaln #(12) e1685(.a(buffered_input), .b(12'b011010010101), .eq(weq1685));
    equaln #(12) e1686(.a(buffered_input), .b(12'b011010010110), .eq(weq1686));
    equaln #(12) e1687(.a(buffered_input), .b(12'b011010010111), .eq(weq1687));
    equaln #(12) e1688(.a(buffered_input), .b(12'b011010011000), .eq(weq1688));
    equaln #(12) e1689(.a(buffered_input), .b(12'b011010011001), .eq(weq1689));
    equaln #(12) e1690(.a(buffered_input), .b(12'b011010011010), .eq(weq1690));
    equaln #(12) e1691(.a(buffered_input), .b(12'b011010011011), .eq(weq1691));
    equaln #(12) e1692(.a(buffered_input), .b(12'b011010011100), .eq(weq1692));
    equaln #(12) e1693(.a(buffered_input), .b(12'b011010011101), .eq(weq1693));
    equaln #(12) e1694(.a(buffered_input), .b(12'b011010011110), .eq(weq1694));
    equaln #(12) e1695(.a(buffered_input), .b(12'b011010011111), .eq(weq1695));
    equaln #(12) e1696(.a(buffered_input), .b(12'b011010100000), .eq(weq1696));
    equaln #(12) e1697(.a(buffered_input), .b(12'b011010100001), .eq(weq1697));
    equaln #(12) e1698(.a(buffered_input), .b(12'b011010100010), .eq(weq1698));
    equaln #(12) e1699(.a(buffered_input), .b(12'b011010100011), .eq(weq1699));
    equaln #(12) e1700(.a(buffered_input), .b(12'b011010100100), .eq(weq1700));
    equaln #(12) e1701(.a(buffered_input), .b(12'b011010100101), .eq(weq1701));
    equaln #(12) e1702(.a(buffered_input), .b(12'b011010100110), .eq(weq1702));
    equaln #(12) e1703(.a(buffered_input), .b(12'b011010100111), .eq(weq1703));
    equaln #(12) e1704(.a(buffered_input), .b(12'b011010101000), .eq(weq1704));
    equaln #(12) e1705(.a(buffered_input), .b(12'b011010101001), .eq(weq1705));
    equaln #(12) e1706(.a(buffered_input), .b(12'b011010101010), .eq(weq1706));
    equaln #(12) e1707(.a(buffered_input), .b(12'b011010101011), .eq(weq1707));
    equaln #(12) e1708(.a(buffered_input), .b(12'b011010101100), .eq(weq1708));
    equaln #(12) e1709(.a(buffered_input), .b(12'b011010101101), .eq(weq1709));
    equaln #(12) e1710(.a(buffered_input), .b(12'b011010101110), .eq(weq1710));
    equaln #(12) e1711(.a(buffered_input), .b(12'b011010101111), .eq(weq1711));
    equaln #(12) e1712(.a(buffered_input), .b(12'b011010110000), .eq(weq1712));
    equaln #(12) e1713(.a(buffered_input), .b(12'b011010110001), .eq(weq1713));
    equaln #(12) e1714(.a(buffered_input), .b(12'b011010110010), .eq(weq1714));
    equaln #(12) e1715(.a(buffered_input), .b(12'b011010110011), .eq(weq1715));
    equaln #(12) e1716(.a(buffered_input), .b(12'b011010110100), .eq(weq1716));
    equaln #(12) e1717(.a(buffered_input), .b(12'b011010110101), .eq(weq1717));
    equaln #(12) e1718(.a(buffered_input), .b(12'b011010110110), .eq(weq1718));
    equaln #(12) e1719(.a(buffered_input), .b(12'b011010110111), .eq(weq1719));
    equaln #(12) e1720(.a(buffered_input), .b(12'b011010111000), .eq(weq1720));
    equaln #(12) e1721(.a(buffered_input), .b(12'b011010111001), .eq(weq1721));
    equaln #(12) e1722(.a(buffered_input), .b(12'b011010111010), .eq(weq1722));
    equaln #(12) e1723(.a(buffered_input), .b(12'b011010111011), .eq(weq1723));
    equaln #(12) e1724(.a(buffered_input), .b(12'b011010111100), .eq(weq1724));
    equaln #(12) e1725(.a(buffered_input), .b(12'b011010111101), .eq(weq1725));
    equaln #(12) e1726(.a(buffered_input), .b(12'b011010111110), .eq(weq1726));
    equaln #(12) e1727(.a(buffered_input), .b(12'b011010111111), .eq(weq1727));
    equaln #(12) e1728(.a(buffered_input), .b(12'b011011000000), .eq(weq1728));
    equaln #(12) e1729(.a(buffered_input), .b(12'b011011000001), .eq(weq1729));
    equaln #(12) e1730(.a(buffered_input), .b(12'b011011000010), .eq(weq1730));
    equaln #(12) e1731(.a(buffered_input), .b(12'b011011000011), .eq(weq1731));
    equaln #(12) e1732(.a(buffered_input), .b(12'b011011000100), .eq(weq1732));
    equaln #(12) e1733(.a(buffered_input), .b(12'b011011000101), .eq(weq1733));
    equaln #(12) e1734(.a(buffered_input), .b(12'b011011000110), .eq(weq1734));
    equaln #(12) e1735(.a(buffered_input), .b(12'b011011000111), .eq(weq1735));
    equaln #(12) e1736(.a(buffered_input), .b(12'b011011001000), .eq(weq1736));
    equaln #(12) e1737(.a(buffered_input), .b(12'b011011001001), .eq(weq1737));
    equaln #(12) e1738(.a(buffered_input), .b(12'b011011001010), .eq(weq1738));
    equaln #(12) e1739(.a(buffered_input), .b(12'b011011001011), .eq(weq1739));
    equaln #(12) e1740(.a(buffered_input), .b(12'b011011001100), .eq(weq1740));
    equaln #(12) e1741(.a(buffered_input), .b(12'b011011001101), .eq(weq1741));
    equaln #(12) e1742(.a(buffered_input), .b(12'b011011001110), .eq(weq1742));
    equaln #(12) e1743(.a(buffered_input), .b(12'b011011001111), .eq(weq1743));
    equaln #(12) e1744(.a(buffered_input), .b(12'b011011010000), .eq(weq1744));
    equaln #(12) e1745(.a(buffered_input), .b(12'b011011010001), .eq(weq1745));
    equaln #(12) e1746(.a(buffered_input), .b(12'b011011010010), .eq(weq1746));
    equaln #(12) e1747(.a(buffered_input), .b(12'b011011010011), .eq(weq1747));
    equaln #(12) e1748(.a(buffered_input), .b(12'b011011010100), .eq(weq1748));
    equaln #(12) e1749(.a(buffered_input), .b(12'b011011010101), .eq(weq1749));
    equaln #(12) e1750(.a(buffered_input), .b(12'b011011010110), .eq(weq1750));
    equaln #(12) e1751(.a(buffered_input), .b(12'b011011010111), .eq(weq1751));
    equaln #(12) e1752(.a(buffered_input), .b(12'b011011011000), .eq(weq1752));
    equaln #(12) e1753(.a(buffered_input), .b(12'b011011011001), .eq(weq1753));
    equaln #(12) e1754(.a(buffered_input), .b(12'b011011011010), .eq(weq1754));
    equaln #(12) e1755(.a(buffered_input), .b(12'b011011011011), .eq(weq1755));
    equaln #(12) e1756(.a(buffered_input), .b(12'b011011011100), .eq(weq1756));
    equaln #(12) e1757(.a(buffered_input), .b(12'b011011011101), .eq(weq1757));
    equaln #(12) e1758(.a(buffered_input), .b(12'b011011011110), .eq(weq1758));
    equaln #(12) e1759(.a(buffered_input), .b(12'b011011011111), .eq(weq1759));
    equaln #(12) e1760(.a(buffered_input), .b(12'b011011100000), .eq(weq1760));
    equaln #(12) e1761(.a(buffered_input), .b(12'b011011100001), .eq(weq1761));
    equaln #(12) e1762(.a(buffered_input), .b(12'b011011100010), .eq(weq1762));
    equaln #(12) e1763(.a(buffered_input), .b(12'b011011100011), .eq(weq1763));
    equaln #(12) e1764(.a(buffered_input), .b(12'b011011100100), .eq(weq1764));
    equaln #(12) e1765(.a(buffered_input), .b(12'b011011100101), .eq(weq1765));
    equaln #(12) e1766(.a(buffered_input), .b(12'b011011100110), .eq(weq1766));
    equaln #(12) e1767(.a(buffered_input), .b(12'b011011100111), .eq(weq1767));
    equaln #(12) e1768(.a(buffered_input), .b(12'b011011101000), .eq(weq1768));
    equaln #(12) e1769(.a(buffered_input), .b(12'b011011101001), .eq(weq1769));
    equaln #(12) e1770(.a(buffered_input), .b(12'b011011101010), .eq(weq1770));
    equaln #(12) e1771(.a(buffered_input), .b(12'b011011101011), .eq(weq1771));
    equaln #(12) e1772(.a(buffered_input), .b(12'b011011101100), .eq(weq1772));
    equaln #(12) e1773(.a(buffered_input), .b(12'b011011101101), .eq(weq1773));
    equaln #(12) e1774(.a(buffered_input), .b(12'b011011101110), .eq(weq1774));
    equaln #(12) e1775(.a(buffered_input), .b(12'b011011101111), .eq(weq1775));
    equaln #(12) e1776(.a(buffered_input), .b(12'b011011110000), .eq(weq1776));
    equaln #(12) e1777(.a(buffered_input), .b(12'b011011110001), .eq(weq1777));
    equaln #(12) e1778(.a(buffered_input), .b(12'b011011110010), .eq(weq1778));
    equaln #(12) e1779(.a(buffered_input), .b(12'b011011110011), .eq(weq1779));
    equaln #(12) e1780(.a(buffered_input), .b(12'b011011110100), .eq(weq1780));
    equaln #(12) e1781(.a(buffered_input), .b(12'b011011110101), .eq(weq1781));
    equaln #(12) e1782(.a(buffered_input), .b(12'b011011110110), .eq(weq1782));
    equaln #(12) e1783(.a(buffered_input), .b(12'b011011110111), .eq(weq1783));
    equaln #(12) e1784(.a(buffered_input), .b(12'b011011111000), .eq(weq1784));
    equaln #(12) e1785(.a(buffered_input), .b(12'b011011111001), .eq(weq1785));
    equaln #(12) e1786(.a(buffered_input), .b(12'b011011111010), .eq(weq1786));
    equaln #(12) e1787(.a(buffered_input), .b(12'b011011111011), .eq(weq1787));
    equaln #(12) e1788(.a(buffered_input), .b(12'b011011111100), .eq(weq1788));
    equaln #(12) e1789(.a(buffered_input), .b(12'b011011111101), .eq(weq1789));
    equaln #(12) e1790(.a(buffered_input), .b(12'b011011111110), .eq(weq1790));
    equaln #(12) e1791(.a(buffered_input), .b(12'b011011111111), .eq(weq1791));
    equaln #(12) e1792(.a(buffered_input), .b(12'b011100000000), .eq(weq1792));
    equaln #(12) e1793(.a(buffered_input), .b(12'b011100000001), .eq(weq1793));
    equaln #(12) e1794(.a(buffered_input), .b(12'b011100000010), .eq(weq1794));
    equaln #(12) e1795(.a(buffered_input), .b(12'b011100000011), .eq(weq1795));
    equaln #(12) e1796(.a(buffered_input), .b(12'b011100000100), .eq(weq1796));
    equaln #(12) e1797(.a(buffered_input), .b(12'b011100000101), .eq(weq1797));
    equaln #(12) e1798(.a(buffered_input), .b(12'b011100000110), .eq(weq1798));
    equaln #(12) e1799(.a(buffered_input), .b(12'b011100000111), .eq(weq1799));
    equaln #(12) e1800(.a(buffered_input), .b(12'b011100001000), .eq(weq1800));
    equaln #(12) e1801(.a(buffered_input), .b(12'b011100001001), .eq(weq1801));
    equaln #(12) e1802(.a(buffered_input), .b(12'b011100001010), .eq(weq1802));
    equaln #(12) e1803(.a(buffered_input), .b(12'b011100001011), .eq(weq1803));
    equaln #(12) e1804(.a(buffered_input), .b(12'b011100001100), .eq(weq1804));
    equaln #(12) e1805(.a(buffered_input), .b(12'b011100001101), .eq(weq1805));
    equaln #(12) e1806(.a(buffered_input), .b(12'b011100001110), .eq(weq1806));
    equaln #(12) e1807(.a(buffered_input), .b(12'b011100001111), .eq(weq1807));
    equaln #(12) e1808(.a(buffered_input), .b(12'b011100010000), .eq(weq1808));
    equaln #(12) e1809(.a(buffered_input), .b(12'b011100010001), .eq(weq1809));
    equaln #(12) e1810(.a(buffered_input), .b(12'b011100010010), .eq(weq1810));
    equaln #(12) e1811(.a(buffered_input), .b(12'b011100010011), .eq(weq1811));
    equaln #(12) e1812(.a(buffered_input), .b(12'b011100010100), .eq(weq1812));
    equaln #(12) e1813(.a(buffered_input), .b(12'b011100010101), .eq(weq1813));
    equaln #(12) e1814(.a(buffered_input), .b(12'b011100010110), .eq(weq1814));
    equaln #(12) e1815(.a(buffered_input), .b(12'b011100010111), .eq(weq1815));
    equaln #(12) e1816(.a(buffered_input), .b(12'b011100011000), .eq(weq1816));
    equaln #(12) e1817(.a(buffered_input), .b(12'b011100011001), .eq(weq1817));
    equaln #(12) e1818(.a(buffered_input), .b(12'b011100011010), .eq(weq1818));
    equaln #(12) e1819(.a(buffered_input), .b(12'b011100011011), .eq(weq1819));
    equaln #(12) e1820(.a(buffered_input), .b(12'b011100011100), .eq(weq1820));
    equaln #(12) e1821(.a(buffered_input), .b(12'b011100011101), .eq(weq1821));
    equaln #(12) e1822(.a(buffered_input), .b(12'b011100011110), .eq(weq1822));
    equaln #(12) e1823(.a(buffered_input), .b(12'b011100011111), .eq(weq1823));
    equaln #(12) e1824(.a(buffered_input), .b(12'b011100100000), .eq(weq1824));
    equaln #(12) e1825(.a(buffered_input), .b(12'b011100100001), .eq(weq1825));
    equaln #(12) e1826(.a(buffered_input), .b(12'b011100100010), .eq(weq1826));
    equaln #(12) e1827(.a(buffered_input), .b(12'b011100100011), .eq(weq1827));
    equaln #(12) e1828(.a(buffered_input), .b(12'b011100100100), .eq(weq1828));
    equaln #(12) e1829(.a(buffered_input), .b(12'b011100100101), .eq(weq1829));
    equaln #(12) e1830(.a(buffered_input), .b(12'b011100100110), .eq(weq1830));
    equaln #(12) e1831(.a(buffered_input), .b(12'b011100100111), .eq(weq1831));
    equaln #(12) e1832(.a(buffered_input), .b(12'b011100101000), .eq(weq1832));
    equaln #(12) e1833(.a(buffered_input), .b(12'b011100101001), .eq(weq1833));
    equaln #(12) e1834(.a(buffered_input), .b(12'b011100101010), .eq(weq1834));
    equaln #(12) e1835(.a(buffered_input), .b(12'b011100101011), .eq(weq1835));
    equaln #(12) e1836(.a(buffered_input), .b(12'b011100101100), .eq(weq1836));
    equaln #(12) e1837(.a(buffered_input), .b(12'b011100101101), .eq(weq1837));
    equaln #(12) e1838(.a(buffered_input), .b(12'b011100101110), .eq(weq1838));
    equaln #(12) e1839(.a(buffered_input), .b(12'b011100101111), .eq(weq1839));
    equaln #(12) e1840(.a(buffered_input), .b(12'b011100110000), .eq(weq1840));
    equaln #(12) e1841(.a(buffered_input), .b(12'b011100110001), .eq(weq1841));
    equaln #(12) e1842(.a(buffered_input), .b(12'b011100110010), .eq(weq1842));
    equaln #(12) e1843(.a(buffered_input), .b(12'b011100110011), .eq(weq1843));
    equaln #(12) e1844(.a(buffered_input), .b(12'b011100110100), .eq(weq1844));
    equaln #(12) e1845(.a(buffered_input), .b(12'b011100110101), .eq(weq1845));
    equaln #(12) e1846(.a(buffered_input), .b(12'b011100110110), .eq(weq1846));
    equaln #(12) e1847(.a(buffered_input), .b(12'b011100110111), .eq(weq1847));
    equaln #(12) e1848(.a(buffered_input), .b(12'b011100111000), .eq(weq1848));
    equaln #(12) e1849(.a(buffered_input), .b(12'b011100111001), .eq(weq1849));
    equaln #(12) e1850(.a(buffered_input), .b(12'b011100111010), .eq(weq1850));
    equaln #(12) e1851(.a(buffered_input), .b(12'b011100111011), .eq(weq1851));
    equaln #(12) e1852(.a(buffered_input), .b(12'b011100111100), .eq(weq1852));
    equaln #(12) e1853(.a(buffered_input), .b(12'b011100111101), .eq(weq1853));
    equaln #(12) e1854(.a(buffered_input), .b(12'b011100111110), .eq(weq1854));
    equaln #(12) e1855(.a(buffered_input), .b(12'b011100111111), .eq(weq1855));
    equaln #(12) e1856(.a(buffered_input), .b(12'b011101000000), .eq(weq1856));
    equaln #(12) e1857(.a(buffered_input), .b(12'b011101000001), .eq(weq1857));
    equaln #(12) e1858(.a(buffered_input), .b(12'b011101000010), .eq(weq1858));
    equaln #(12) e1859(.a(buffered_input), .b(12'b011101000011), .eq(weq1859));
    equaln #(12) e1860(.a(buffered_input), .b(12'b011101000100), .eq(weq1860));
    equaln #(12) e1861(.a(buffered_input), .b(12'b011101000101), .eq(weq1861));
    equaln #(12) e1862(.a(buffered_input), .b(12'b011101000110), .eq(weq1862));
    equaln #(12) e1863(.a(buffered_input), .b(12'b011101000111), .eq(weq1863));
    equaln #(12) e1864(.a(buffered_input), .b(12'b011101001000), .eq(weq1864));
    equaln #(12) e1865(.a(buffered_input), .b(12'b011101001001), .eq(weq1865));
    equaln #(12) e1866(.a(buffered_input), .b(12'b011101001010), .eq(weq1866));
    equaln #(12) e1867(.a(buffered_input), .b(12'b011101001011), .eq(weq1867));
    equaln #(12) e1868(.a(buffered_input), .b(12'b011101001100), .eq(weq1868));
    equaln #(12) e1869(.a(buffered_input), .b(12'b011101001101), .eq(weq1869));
    equaln #(12) e1870(.a(buffered_input), .b(12'b011101001110), .eq(weq1870));
    equaln #(12) e1871(.a(buffered_input), .b(12'b011101001111), .eq(weq1871));
    equaln #(12) e1872(.a(buffered_input), .b(12'b011101010000), .eq(weq1872));
    equaln #(12) e1873(.a(buffered_input), .b(12'b011101010001), .eq(weq1873));
    equaln #(12) e1874(.a(buffered_input), .b(12'b011101010010), .eq(weq1874));
    equaln #(12) e1875(.a(buffered_input), .b(12'b011101010011), .eq(weq1875));
    equaln #(12) e1876(.a(buffered_input), .b(12'b011101010100), .eq(weq1876));
    equaln #(12) e1877(.a(buffered_input), .b(12'b011101010101), .eq(weq1877));
    equaln #(12) e1878(.a(buffered_input), .b(12'b011101010110), .eq(weq1878));
    equaln #(12) e1879(.a(buffered_input), .b(12'b011101010111), .eq(weq1879));
    equaln #(12) e1880(.a(buffered_input), .b(12'b011101011000), .eq(weq1880));
    equaln #(12) e1881(.a(buffered_input), .b(12'b011101011001), .eq(weq1881));
    equaln #(12) e1882(.a(buffered_input), .b(12'b011101011010), .eq(weq1882));
    equaln #(12) e1883(.a(buffered_input), .b(12'b011101011011), .eq(weq1883));
    equaln #(12) e1884(.a(buffered_input), .b(12'b011101011100), .eq(weq1884));
    equaln #(12) e1885(.a(buffered_input), .b(12'b011101011101), .eq(weq1885));
    equaln #(12) e1886(.a(buffered_input), .b(12'b011101011110), .eq(weq1886));
    equaln #(12) e1887(.a(buffered_input), .b(12'b011101011111), .eq(weq1887));
    equaln #(12) e1888(.a(buffered_input), .b(12'b011101100000), .eq(weq1888));
    equaln #(12) e1889(.a(buffered_input), .b(12'b011101100001), .eq(weq1889));
    equaln #(12) e1890(.a(buffered_input), .b(12'b011101100010), .eq(weq1890));
    equaln #(12) e1891(.a(buffered_input), .b(12'b011101100011), .eq(weq1891));
    equaln #(12) e1892(.a(buffered_input), .b(12'b011101100100), .eq(weq1892));
    equaln #(12) e1893(.a(buffered_input), .b(12'b011101100101), .eq(weq1893));
    equaln #(12) e1894(.a(buffered_input), .b(12'b011101100110), .eq(weq1894));
    equaln #(12) e1895(.a(buffered_input), .b(12'b011101100111), .eq(weq1895));
    equaln #(12) e1896(.a(buffered_input), .b(12'b011101101000), .eq(weq1896));
    equaln #(12) e1897(.a(buffered_input), .b(12'b011101101001), .eq(weq1897));
    equaln #(12) e1898(.a(buffered_input), .b(12'b011101101010), .eq(weq1898));
    equaln #(12) e1899(.a(buffered_input), .b(12'b011101101011), .eq(weq1899));
    equaln #(12) e1900(.a(buffered_input), .b(12'b011101101100), .eq(weq1900));
    equaln #(12) e1901(.a(buffered_input), .b(12'b011101101101), .eq(weq1901));
    equaln #(12) e1902(.a(buffered_input), .b(12'b011101101110), .eq(weq1902));
    equaln #(12) e1903(.a(buffered_input), .b(12'b011101101111), .eq(weq1903));
    equaln #(12) e1904(.a(buffered_input), .b(12'b011101110000), .eq(weq1904));
    equaln #(12) e1905(.a(buffered_input), .b(12'b011101110001), .eq(weq1905));
    equaln #(12) e1906(.a(buffered_input), .b(12'b011101110010), .eq(weq1906));
    equaln #(12) e1907(.a(buffered_input), .b(12'b011101110011), .eq(weq1907));
    equaln #(12) e1908(.a(buffered_input), .b(12'b011101110100), .eq(weq1908));
    equaln #(12) e1909(.a(buffered_input), .b(12'b011101110101), .eq(weq1909));
    equaln #(12) e1910(.a(buffered_input), .b(12'b011101110110), .eq(weq1910));
    equaln #(12) e1911(.a(buffered_input), .b(12'b011101110111), .eq(weq1911));
    equaln #(12) e1912(.a(buffered_input), .b(12'b011101111000), .eq(weq1912));
    equaln #(12) e1913(.a(buffered_input), .b(12'b011101111001), .eq(weq1913));
    equaln #(12) e1914(.a(buffered_input), .b(12'b011101111010), .eq(weq1914));
    equaln #(12) e1915(.a(buffered_input), .b(12'b011101111011), .eq(weq1915));
    equaln #(12) e1916(.a(buffered_input), .b(12'b011101111100), .eq(weq1916));
    equaln #(12) e1917(.a(buffered_input), .b(12'b011101111101), .eq(weq1917));
    equaln #(12) e1918(.a(buffered_input), .b(12'b011101111110), .eq(weq1918));
    equaln #(12) e1919(.a(buffered_input), .b(12'b011101111111), .eq(weq1919));
    equaln #(12) e1920(.a(buffered_input), .b(12'b011110000000), .eq(weq1920));
    equaln #(12) e1921(.a(buffered_input), .b(12'b011110000001), .eq(weq1921));
    equaln #(12) e1922(.a(buffered_input), .b(12'b011110000010), .eq(weq1922));
    equaln #(12) e1923(.a(buffered_input), .b(12'b011110000011), .eq(weq1923));
    equaln #(12) e1924(.a(buffered_input), .b(12'b011110000100), .eq(weq1924));
    equaln #(12) e1925(.a(buffered_input), .b(12'b011110000101), .eq(weq1925));
    equaln #(12) e1926(.a(buffered_input), .b(12'b011110000110), .eq(weq1926));
    equaln #(12) e1927(.a(buffered_input), .b(12'b011110000111), .eq(weq1927));
    equaln #(12) e1928(.a(buffered_input), .b(12'b011110001000), .eq(weq1928));
    equaln #(12) e1929(.a(buffered_input), .b(12'b011110001001), .eq(weq1929));
    equaln #(12) e1930(.a(buffered_input), .b(12'b011110001010), .eq(weq1930));
    equaln #(12) e1931(.a(buffered_input), .b(12'b011110001011), .eq(weq1931));
    equaln #(12) e1932(.a(buffered_input), .b(12'b011110001100), .eq(weq1932));
    equaln #(12) e1933(.a(buffered_input), .b(12'b011110001101), .eq(weq1933));
    equaln #(12) e1934(.a(buffered_input), .b(12'b011110001110), .eq(weq1934));
    equaln #(12) e1935(.a(buffered_input), .b(12'b011110001111), .eq(weq1935));
    equaln #(12) e1936(.a(buffered_input), .b(12'b011110010000), .eq(weq1936));
    equaln #(12) e1937(.a(buffered_input), .b(12'b011110010001), .eq(weq1937));
    equaln #(12) e1938(.a(buffered_input), .b(12'b011110010010), .eq(weq1938));
    equaln #(12) e1939(.a(buffered_input), .b(12'b011110010011), .eq(weq1939));
    equaln #(12) e1940(.a(buffered_input), .b(12'b011110010100), .eq(weq1940));
    equaln #(12) e1941(.a(buffered_input), .b(12'b011110010101), .eq(weq1941));
    equaln #(12) e1942(.a(buffered_input), .b(12'b011110010110), .eq(weq1942));
    equaln #(12) e1943(.a(buffered_input), .b(12'b011110010111), .eq(weq1943));
    equaln #(12) e1944(.a(buffered_input), .b(12'b011110011000), .eq(weq1944));
    equaln #(12) e1945(.a(buffered_input), .b(12'b011110011001), .eq(weq1945));
    equaln #(12) e1946(.a(buffered_input), .b(12'b011110011010), .eq(weq1946));
    equaln #(12) e1947(.a(buffered_input), .b(12'b011110011011), .eq(weq1947));
    equaln #(12) e1948(.a(buffered_input), .b(12'b011110011100), .eq(weq1948));
    equaln #(12) e1949(.a(buffered_input), .b(12'b011110011101), .eq(weq1949));
    equaln #(12) e1950(.a(buffered_input), .b(12'b011110011110), .eq(weq1950));
    equaln #(12) e1951(.a(buffered_input), .b(12'b011110011111), .eq(weq1951));
    equaln #(12) e1952(.a(buffered_input), .b(12'b011110100000), .eq(weq1952));
    equaln #(12) e1953(.a(buffered_input), .b(12'b011110100001), .eq(weq1953));
    equaln #(12) e1954(.a(buffered_input), .b(12'b011110100010), .eq(weq1954));
    equaln #(12) e1955(.a(buffered_input), .b(12'b011110100011), .eq(weq1955));
    equaln #(12) e1956(.a(buffered_input), .b(12'b011110100100), .eq(weq1956));
    equaln #(12) e1957(.a(buffered_input), .b(12'b011110100101), .eq(weq1957));
    equaln #(12) e1958(.a(buffered_input), .b(12'b011110100110), .eq(weq1958));
    equaln #(12) e1959(.a(buffered_input), .b(12'b011110100111), .eq(weq1959));
    equaln #(12) e1960(.a(buffered_input), .b(12'b011110101000), .eq(weq1960));
    equaln #(12) e1961(.a(buffered_input), .b(12'b011110101001), .eq(weq1961));
    equaln #(12) e1962(.a(buffered_input), .b(12'b011110101010), .eq(weq1962));
    equaln #(12) e1963(.a(buffered_input), .b(12'b011110101011), .eq(weq1963));
    equaln #(12) e1964(.a(buffered_input), .b(12'b011110101100), .eq(weq1964));
    equaln #(12) e1965(.a(buffered_input), .b(12'b011110101101), .eq(weq1965));
    equaln #(12) e1966(.a(buffered_input), .b(12'b011110101110), .eq(weq1966));
    equaln #(12) e1967(.a(buffered_input), .b(12'b011110101111), .eq(weq1967));
    equaln #(12) e1968(.a(buffered_input), .b(12'b011110110000), .eq(weq1968));
    equaln #(12) e1969(.a(buffered_input), .b(12'b011110110001), .eq(weq1969));
    equaln #(12) e1970(.a(buffered_input), .b(12'b011110110010), .eq(weq1970));
    equaln #(12) e1971(.a(buffered_input), .b(12'b011110110011), .eq(weq1971));
    equaln #(12) e1972(.a(buffered_input), .b(12'b011110110100), .eq(weq1972));
    equaln #(12) e1973(.a(buffered_input), .b(12'b011110110101), .eq(weq1973));
    equaln #(12) e1974(.a(buffered_input), .b(12'b011110110110), .eq(weq1974));
    equaln #(12) e1975(.a(buffered_input), .b(12'b011110110111), .eq(weq1975));
    equaln #(12) e1976(.a(buffered_input), .b(12'b011110111000), .eq(weq1976));
    equaln #(12) e1977(.a(buffered_input), .b(12'b011110111001), .eq(weq1977));
    equaln #(12) e1978(.a(buffered_input), .b(12'b011110111010), .eq(weq1978));
    equaln #(12) e1979(.a(buffered_input), .b(12'b011110111011), .eq(weq1979));
    equaln #(12) e1980(.a(buffered_input), .b(12'b011110111100), .eq(weq1980));
    equaln #(12) e1981(.a(buffered_input), .b(12'b011110111101), .eq(weq1981));
    equaln #(12) e1982(.a(buffered_input), .b(12'b011110111110), .eq(weq1982));
    equaln #(12) e1983(.a(buffered_input), .b(12'b011110111111), .eq(weq1983));
    equaln #(12) e1984(.a(buffered_input), .b(12'b011111000000), .eq(weq1984));
    equaln #(12) e1985(.a(buffered_input), .b(12'b011111000001), .eq(weq1985));
    equaln #(12) e1986(.a(buffered_input), .b(12'b011111000010), .eq(weq1986));
    equaln #(12) e1987(.a(buffered_input), .b(12'b011111000011), .eq(weq1987));
    equaln #(12) e1988(.a(buffered_input), .b(12'b011111000100), .eq(weq1988));
    equaln #(12) e1989(.a(buffered_input), .b(12'b011111000101), .eq(weq1989));
    equaln #(12) e1990(.a(buffered_input), .b(12'b011111000110), .eq(weq1990));
    equaln #(12) e1991(.a(buffered_input), .b(12'b011111000111), .eq(weq1991));
    equaln #(12) e1992(.a(buffered_input), .b(12'b011111001000), .eq(weq1992));
    equaln #(12) e1993(.a(buffered_input), .b(12'b011111001001), .eq(weq1993));
    equaln #(12) e1994(.a(buffered_input), .b(12'b011111001010), .eq(weq1994));
    equaln #(12) e1995(.a(buffered_input), .b(12'b011111001011), .eq(weq1995));
    equaln #(12) e1996(.a(buffered_input), .b(12'b011111001100), .eq(weq1996));
    equaln #(12) e1997(.a(buffered_input), .b(12'b011111001101), .eq(weq1997));
    equaln #(12) e1998(.a(buffered_input), .b(12'b011111001110), .eq(weq1998));
    equaln #(12) e1999(.a(buffered_input), .b(12'b011111001111), .eq(weq1999));
    equaln #(12) e2000(.a(buffered_input), .b(12'b011111010000), .eq(weq2000));
    equaln #(12) e2001(.a(buffered_input), .b(12'b011111010001), .eq(weq2001));
    equaln #(12) e2002(.a(buffered_input), .b(12'b011111010010), .eq(weq2002));
    equaln #(12) e2003(.a(buffered_input), .b(12'b011111010011), .eq(weq2003));
    equaln #(12) e2004(.a(buffered_input), .b(12'b011111010100), .eq(weq2004));
    equaln #(12) e2005(.a(buffered_input), .b(12'b011111010101), .eq(weq2005));
    equaln #(12) e2006(.a(buffered_input), .b(12'b011111010110), .eq(weq2006));
    equaln #(12) e2007(.a(buffered_input), .b(12'b011111010111), .eq(weq2007));
    equaln #(12) e2008(.a(buffered_input), .b(12'b011111011000), .eq(weq2008));
    equaln #(12) e2009(.a(buffered_input), .b(12'b011111011001), .eq(weq2009));
    equaln #(12) e2010(.a(buffered_input), .b(12'b011111011010), .eq(weq2010));
    equaln #(12) e2011(.a(buffered_input), .b(12'b011111011011), .eq(weq2011));
    equaln #(12) e2012(.a(buffered_input), .b(12'b011111011100), .eq(weq2012));
    equaln #(12) e2013(.a(buffered_input), .b(12'b011111011101), .eq(weq2013));
    equaln #(12) e2014(.a(buffered_input), .b(12'b011111011110), .eq(weq2014));
    equaln #(12) e2015(.a(buffered_input), .b(12'b011111011111), .eq(weq2015));
    equaln #(12) e2016(.a(buffered_input), .b(12'b011111100000), .eq(weq2016));
    equaln #(12) e2017(.a(buffered_input), .b(12'b011111100001), .eq(weq2017));
    equaln #(12) e2018(.a(buffered_input), .b(12'b011111100010), .eq(weq2018));
    equaln #(12) e2019(.a(buffered_input), .b(12'b011111100011), .eq(weq2019));
    equaln #(12) e2020(.a(buffered_input), .b(12'b011111100100), .eq(weq2020));
    equaln #(12) e2021(.a(buffered_input), .b(12'b011111100101), .eq(weq2021));
    equaln #(12) e2022(.a(buffered_input), .b(12'b011111100110), .eq(weq2022));
    equaln #(12) e2023(.a(buffered_input), .b(12'b011111100111), .eq(weq2023));
    equaln #(12) e2024(.a(buffered_input), .b(12'b011111101000), .eq(weq2024));
    equaln #(12) e2025(.a(buffered_input), .b(12'b011111101001), .eq(weq2025));
    equaln #(12) e2026(.a(buffered_input), .b(12'b011111101010), .eq(weq2026));
    equaln #(12) e2027(.a(buffered_input), .b(12'b011111101011), .eq(weq2027));
    equaln #(12) e2028(.a(buffered_input), .b(12'b011111101100), .eq(weq2028));
    equaln #(12) e2029(.a(buffered_input), .b(12'b011111101101), .eq(weq2029));
    equaln #(12) e2030(.a(buffered_input), .b(12'b011111101110), .eq(weq2030));
    equaln #(12) e2031(.a(buffered_input), .b(12'b011111101111), .eq(weq2031));
    equaln #(12) e2032(.a(buffered_input), .b(12'b011111110000), .eq(weq2032));
    equaln #(12) e2033(.a(buffered_input), .b(12'b011111110001), .eq(weq2033));
    equaln #(12) e2034(.a(buffered_input), .b(12'b011111110010), .eq(weq2034));
    equaln #(12) e2035(.a(buffered_input), .b(12'b011111110011), .eq(weq2035));
    equaln #(12) e2036(.a(buffered_input), .b(12'b011111110100), .eq(weq2036));
    equaln #(12) e2037(.a(buffered_input), .b(12'b011111110101), .eq(weq2037));
    equaln #(12) e2038(.a(buffered_input), .b(12'b011111110110), .eq(weq2038));
    equaln #(12) e2039(.a(buffered_input), .b(12'b011111110111), .eq(weq2039));
    equaln #(12) e2040(.a(buffered_input), .b(12'b011111111000), .eq(weq2040));
    equaln #(12) e2041(.a(buffered_input), .b(12'b011111111001), .eq(weq2041));
    equaln #(12) e2042(.a(buffered_input), .b(12'b011111111010), .eq(weq2042));
    equaln #(12) e2043(.a(buffered_input), .b(12'b011111111011), .eq(weq2043));
    equaln #(12) e2044(.a(buffered_input), .b(12'b011111111100), .eq(weq2044));
    equaln #(12) e2045(.a(buffered_input), .b(12'b011111111101), .eq(weq2045));
    equaln #(12) e2046(.a(buffered_input), .b(12'b011111111110), .eq(weq2046));
    equaln #(12) e2047(.a(buffered_input), .b(12'b011111111111), .eq(weq2047));
    equaln #(12) e2048(.a(buffered_input), .b(12'b100000000000), .eq(weq2048));
    equaln #(12) e2049(.a(buffered_input), .b(12'b100000000001), .eq(weq2049));
    equaln #(12) e2050(.a(buffered_input), .b(12'b100000000010), .eq(weq2050));
    equaln #(12) e2051(.a(buffered_input), .b(12'b100000000011), .eq(weq2051));
    equaln #(12) e2052(.a(buffered_input), .b(12'b100000000100), .eq(weq2052));
    equaln #(12) e2053(.a(buffered_input), .b(12'b100000000101), .eq(weq2053));
    equaln #(12) e2054(.a(buffered_input), .b(12'b100000000110), .eq(weq2054));
    equaln #(12) e2055(.a(buffered_input), .b(12'b100000000111), .eq(weq2055));
    equaln #(12) e2056(.a(buffered_input), .b(12'b100000001000), .eq(weq2056));
    equaln #(12) e2057(.a(buffered_input), .b(12'b100000001001), .eq(weq2057));
    equaln #(12) e2058(.a(buffered_input), .b(12'b100000001010), .eq(weq2058));
    equaln #(12) e2059(.a(buffered_input), .b(12'b100000001011), .eq(weq2059));
    equaln #(12) e2060(.a(buffered_input), .b(12'b100000001100), .eq(weq2060));
    equaln #(12) e2061(.a(buffered_input), .b(12'b100000001101), .eq(weq2061));
    equaln #(12) e2062(.a(buffered_input), .b(12'b100000001110), .eq(weq2062));
    equaln #(12) e2063(.a(buffered_input), .b(12'b100000001111), .eq(weq2063));
    equaln #(12) e2064(.a(buffered_input), .b(12'b100000010000), .eq(weq2064));
    equaln #(12) e2065(.a(buffered_input), .b(12'b100000010001), .eq(weq2065));
    equaln #(12) e2066(.a(buffered_input), .b(12'b100000010010), .eq(weq2066));
    equaln #(12) e2067(.a(buffered_input), .b(12'b100000010011), .eq(weq2067));
    equaln #(12) e2068(.a(buffered_input), .b(12'b100000010100), .eq(weq2068));
    equaln #(12) e2069(.a(buffered_input), .b(12'b100000010101), .eq(weq2069));
    equaln #(12) e2070(.a(buffered_input), .b(12'b100000010110), .eq(weq2070));
    equaln #(12) e2071(.a(buffered_input), .b(12'b100000010111), .eq(weq2071));
    equaln #(12) e2072(.a(buffered_input), .b(12'b100000011000), .eq(weq2072));
    equaln #(12) e2073(.a(buffered_input), .b(12'b100000011001), .eq(weq2073));
    equaln #(12) e2074(.a(buffered_input), .b(12'b100000011010), .eq(weq2074));
    equaln #(12) e2075(.a(buffered_input), .b(12'b100000011011), .eq(weq2075));
    equaln #(12) e2076(.a(buffered_input), .b(12'b100000011100), .eq(weq2076));
    equaln #(12) e2077(.a(buffered_input), .b(12'b100000011101), .eq(weq2077));
    equaln #(12) e2078(.a(buffered_input), .b(12'b100000011110), .eq(weq2078));
    equaln #(12) e2079(.a(buffered_input), .b(12'b100000011111), .eq(weq2079));
    equaln #(12) e2080(.a(buffered_input), .b(12'b100000100000), .eq(weq2080));
    equaln #(12) e2081(.a(buffered_input), .b(12'b100000100001), .eq(weq2081));
    equaln #(12) e2082(.a(buffered_input), .b(12'b100000100010), .eq(weq2082));
    equaln #(12) e2083(.a(buffered_input), .b(12'b100000100011), .eq(weq2083));
    equaln #(12) e2084(.a(buffered_input), .b(12'b100000100100), .eq(weq2084));
    equaln #(12) e2085(.a(buffered_input), .b(12'b100000100101), .eq(weq2085));
    equaln #(12) e2086(.a(buffered_input), .b(12'b100000100110), .eq(weq2086));
    equaln #(12) e2087(.a(buffered_input), .b(12'b100000100111), .eq(weq2087));
    equaln #(12) e2088(.a(buffered_input), .b(12'b100000101000), .eq(weq2088));
    equaln #(12) e2089(.a(buffered_input), .b(12'b100000101001), .eq(weq2089));
    equaln #(12) e2090(.a(buffered_input), .b(12'b100000101010), .eq(weq2090));
    equaln #(12) e2091(.a(buffered_input), .b(12'b100000101011), .eq(weq2091));
    equaln #(12) e2092(.a(buffered_input), .b(12'b100000101100), .eq(weq2092));
    equaln #(12) e2093(.a(buffered_input), .b(12'b100000101101), .eq(weq2093));
    equaln #(12) e2094(.a(buffered_input), .b(12'b100000101110), .eq(weq2094));
    equaln #(12) e2095(.a(buffered_input), .b(12'b100000101111), .eq(weq2095));
    equaln #(12) e2096(.a(buffered_input), .b(12'b100000110000), .eq(weq2096));
    equaln #(12) e2097(.a(buffered_input), .b(12'b100000110001), .eq(weq2097));
    equaln #(12) e2098(.a(buffered_input), .b(12'b100000110010), .eq(weq2098));
    equaln #(12) e2099(.a(buffered_input), .b(12'b100000110011), .eq(weq2099));
    equaln #(12) e2100(.a(buffered_input), .b(12'b100000110100), .eq(weq2100));
    equaln #(12) e2101(.a(buffered_input), .b(12'b100000110101), .eq(weq2101));
    equaln #(12) e2102(.a(buffered_input), .b(12'b100000110110), .eq(weq2102));
    equaln #(12) e2103(.a(buffered_input), .b(12'b100000110111), .eq(weq2103));
    equaln #(12) e2104(.a(buffered_input), .b(12'b100000111000), .eq(weq2104));
    equaln #(12) e2105(.a(buffered_input), .b(12'b100000111001), .eq(weq2105));
    equaln #(12) e2106(.a(buffered_input), .b(12'b100000111010), .eq(weq2106));
    equaln #(12) e2107(.a(buffered_input), .b(12'b100000111011), .eq(weq2107));
    equaln #(12) e2108(.a(buffered_input), .b(12'b100000111100), .eq(weq2108));
    equaln #(12) e2109(.a(buffered_input), .b(12'b100000111101), .eq(weq2109));
    equaln #(12) e2110(.a(buffered_input), .b(12'b100000111110), .eq(weq2110));
    equaln #(12) e2111(.a(buffered_input), .b(12'b100000111111), .eq(weq2111));
    equaln #(12) e2112(.a(buffered_input), .b(12'b100001000000), .eq(weq2112));
    equaln #(12) e2113(.a(buffered_input), .b(12'b100001000001), .eq(weq2113));
    equaln #(12) e2114(.a(buffered_input), .b(12'b100001000010), .eq(weq2114));
    equaln #(12) e2115(.a(buffered_input), .b(12'b100001000011), .eq(weq2115));
    equaln #(12) e2116(.a(buffered_input), .b(12'b100001000100), .eq(weq2116));
    equaln #(12) e2117(.a(buffered_input), .b(12'b100001000101), .eq(weq2117));
    equaln #(12) e2118(.a(buffered_input), .b(12'b100001000110), .eq(weq2118));
    equaln #(12) e2119(.a(buffered_input), .b(12'b100001000111), .eq(weq2119));
    equaln #(12) e2120(.a(buffered_input), .b(12'b100001001000), .eq(weq2120));
    equaln #(12) e2121(.a(buffered_input), .b(12'b100001001001), .eq(weq2121));
    equaln #(12) e2122(.a(buffered_input), .b(12'b100001001010), .eq(weq2122));
    equaln #(12) e2123(.a(buffered_input), .b(12'b100001001011), .eq(weq2123));
    equaln #(12) e2124(.a(buffered_input), .b(12'b100001001100), .eq(weq2124));
    equaln #(12) e2125(.a(buffered_input), .b(12'b100001001101), .eq(weq2125));
    equaln #(12) e2126(.a(buffered_input), .b(12'b100001001110), .eq(weq2126));
    equaln #(12) e2127(.a(buffered_input), .b(12'b100001001111), .eq(weq2127));
    equaln #(12) e2128(.a(buffered_input), .b(12'b100001010000), .eq(weq2128));
    equaln #(12) e2129(.a(buffered_input), .b(12'b100001010001), .eq(weq2129));
    equaln #(12) e2130(.a(buffered_input), .b(12'b100001010010), .eq(weq2130));
    equaln #(12) e2131(.a(buffered_input), .b(12'b100001010011), .eq(weq2131));
    equaln #(12) e2132(.a(buffered_input), .b(12'b100001010100), .eq(weq2132));
    equaln #(12) e2133(.a(buffered_input), .b(12'b100001010101), .eq(weq2133));
    equaln #(12) e2134(.a(buffered_input), .b(12'b100001010110), .eq(weq2134));
    equaln #(12) e2135(.a(buffered_input), .b(12'b100001010111), .eq(weq2135));
    equaln #(12) e2136(.a(buffered_input), .b(12'b100001011000), .eq(weq2136));
    equaln #(12) e2137(.a(buffered_input), .b(12'b100001011001), .eq(weq2137));
    equaln #(12) e2138(.a(buffered_input), .b(12'b100001011010), .eq(weq2138));
    equaln #(12) e2139(.a(buffered_input), .b(12'b100001011011), .eq(weq2139));
    equaln #(12) e2140(.a(buffered_input), .b(12'b100001011100), .eq(weq2140));
    equaln #(12) e2141(.a(buffered_input), .b(12'b100001011101), .eq(weq2141));
    equaln #(12) e2142(.a(buffered_input), .b(12'b100001011110), .eq(weq2142));
    equaln #(12) e2143(.a(buffered_input), .b(12'b100001011111), .eq(weq2143));
    equaln #(12) e2144(.a(buffered_input), .b(12'b100001100000), .eq(weq2144));
    equaln #(12) e2145(.a(buffered_input), .b(12'b100001100001), .eq(weq2145));
    equaln #(12) e2146(.a(buffered_input), .b(12'b100001100010), .eq(weq2146));
    equaln #(12) e2147(.a(buffered_input), .b(12'b100001100011), .eq(weq2147));
    equaln #(12) e2148(.a(buffered_input), .b(12'b100001100100), .eq(weq2148));
    equaln #(12) e2149(.a(buffered_input), .b(12'b100001100101), .eq(weq2149));
    equaln #(12) e2150(.a(buffered_input), .b(12'b100001100110), .eq(weq2150));
    equaln #(12) e2151(.a(buffered_input), .b(12'b100001100111), .eq(weq2151));
    equaln #(12) e2152(.a(buffered_input), .b(12'b100001101000), .eq(weq2152));
    equaln #(12) e2153(.a(buffered_input), .b(12'b100001101001), .eq(weq2153));
    equaln #(12) e2154(.a(buffered_input), .b(12'b100001101010), .eq(weq2154));
    equaln #(12) e2155(.a(buffered_input), .b(12'b100001101011), .eq(weq2155));
    equaln #(12) e2156(.a(buffered_input), .b(12'b100001101100), .eq(weq2156));
    equaln #(12) e2157(.a(buffered_input), .b(12'b100001101101), .eq(weq2157));
    equaln #(12) e2158(.a(buffered_input), .b(12'b100001101110), .eq(weq2158));
    equaln #(12) e2159(.a(buffered_input), .b(12'b100001101111), .eq(weq2159));
    equaln #(12) e2160(.a(buffered_input), .b(12'b100001110000), .eq(weq2160));
    equaln #(12) e2161(.a(buffered_input), .b(12'b100001110001), .eq(weq2161));
    equaln #(12) e2162(.a(buffered_input), .b(12'b100001110010), .eq(weq2162));
    equaln #(12) e2163(.a(buffered_input), .b(12'b100001110011), .eq(weq2163));
    equaln #(12) e2164(.a(buffered_input), .b(12'b100001110100), .eq(weq2164));
    equaln #(12) e2165(.a(buffered_input), .b(12'b100001110101), .eq(weq2165));
    equaln #(12) e2166(.a(buffered_input), .b(12'b100001110110), .eq(weq2166));
    equaln #(12) e2167(.a(buffered_input), .b(12'b100001110111), .eq(weq2167));
    equaln #(12) e2168(.a(buffered_input), .b(12'b100001111000), .eq(weq2168));
    equaln #(12) e2169(.a(buffered_input), .b(12'b100001111001), .eq(weq2169));
    equaln #(12) e2170(.a(buffered_input), .b(12'b100001111010), .eq(weq2170));
    equaln #(12) e2171(.a(buffered_input), .b(12'b100001111011), .eq(weq2171));
    equaln #(12) e2172(.a(buffered_input), .b(12'b100001111100), .eq(weq2172));
    equaln #(12) e2173(.a(buffered_input), .b(12'b100001111101), .eq(weq2173));
    equaln #(12) e2174(.a(buffered_input), .b(12'b100001111110), .eq(weq2174));
    equaln #(12) e2175(.a(buffered_input), .b(12'b100001111111), .eq(weq2175));
    equaln #(12) e2176(.a(buffered_input), .b(12'b100010000000), .eq(weq2176));
    equaln #(12) e2177(.a(buffered_input), .b(12'b100010000001), .eq(weq2177));
    equaln #(12) e2178(.a(buffered_input), .b(12'b100010000010), .eq(weq2178));
    equaln #(12) e2179(.a(buffered_input), .b(12'b100010000011), .eq(weq2179));
    equaln #(12) e2180(.a(buffered_input), .b(12'b100010000100), .eq(weq2180));
    equaln #(12) e2181(.a(buffered_input), .b(12'b100010000101), .eq(weq2181));
    equaln #(12) e2182(.a(buffered_input), .b(12'b100010000110), .eq(weq2182));
    equaln #(12) e2183(.a(buffered_input), .b(12'b100010000111), .eq(weq2183));
    equaln #(12) e2184(.a(buffered_input), .b(12'b100010001000), .eq(weq2184));
    equaln #(12) e2185(.a(buffered_input), .b(12'b100010001001), .eq(weq2185));
    equaln #(12) e2186(.a(buffered_input), .b(12'b100010001010), .eq(weq2186));
    equaln #(12) e2187(.a(buffered_input), .b(12'b100010001011), .eq(weq2187));
    equaln #(12) e2188(.a(buffered_input), .b(12'b100010001100), .eq(weq2188));
    equaln #(12) e2189(.a(buffered_input), .b(12'b100010001101), .eq(weq2189));
    equaln #(12) e2190(.a(buffered_input), .b(12'b100010001110), .eq(weq2190));
    equaln #(12) e2191(.a(buffered_input), .b(12'b100010001111), .eq(weq2191));
    equaln #(12) e2192(.a(buffered_input), .b(12'b100010010000), .eq(weq2192));
    equaln #(12) e2193(.a(buffered_input), .b(12'b100010010001), .eq(weq2193));
    equaln #(12) e2194(.a(buffered_input), .b(12'b100010010010), .eq(weq2194));
    equaln #(12) e2195(.a(buffered_input), .b(12'b100010010011), .eq(weq2195));
    equaln #(12) e2196(.a(buffered_input), .b(12'b100010010100), .eq(weq2196));
    equaln #(12) e2197(.a(buffered_input), .b(12'b100010010101), .eq(weq2197));
    equaln #(12) e2198(.a(buffered_input), .b(12'b100010010110), .eq(weq2198));
    equaln #(12) e2199(.a(buffered_input), .b(12'b100010010111), .eq(weq2199));
    equaln #(12) e2200(.a(buffered_input), .b(12'b100010011000), .eq(weq2200));
    equaln #(12) e2201(.a(buffered_input), .b(12'b100010011001), .eq(weq2201));
    equaln #(12) e2202(.a(buffered_input), .b(12'b100010011010), .eq(weq2202));
    equaln #(12) e2203(.a(buffered_input), .b(12'b100010011011), .eq(weq2203));
    equaln #(12) e2204(.a(buffered_input), .b(12'b100010011100), .eq(weq2204));
    equaln #(12) e2205(.a(buffered_input), .b(12'b100010011101), .eq(weq2205));
    equaln #(12) e2206(.a(buffered_input), .b(12'b100010011110), .eq(weq2206));
    equaln #(12) e2207(.a(buffered_input), .b(12'b100010011111), .eq(weq2207));
    equaln #(12) e2208(.a(buffered_input), .b(12'b100010100000), .eq(weq2208));
    equaln #(12) e2209(.a(buffered_input), .b(12'b100010100001), .eq(weq2209));
    equaln #(12) e2210(.a(buffered_input), .b(12'b100010100010), .eq(weq2210));
    equaln #(12) e2211(.a(buffered_input), .b(12'b100010100011), .eq(weq2211));
    equaln #(12) e2212(.a(buffered_input), .b(12'b100010100100), .eq(weq2212));
    equaln #(12) e2213(.a(buffered_input), .b(12'b100010100101), .eq(weq2213));
    equaln #(12) e2214(.a(buffered_input), .b(12'b100010100110), .eq(weq2214));
    equaln #(12) e2215(.a(buffered_input), .b(12'b100010100111), .eq(weq2215));
    equaln #(12) e2216(.a(buffered_input), .b(12'b100010101000), .eq(weq2216));
    equaln #(12) e2217(.a(buffered_input), .b(12'b100010101001), .eq(weq2217));
    equaln #(12) e2218(.a(buffered_input), .b(12'b100010101010), .eq(weq2218));
    equaln #(12) e2219(.a(buffered_input), .b(12'b100010101011), .eq(weq2219));
    equaln #(12) e2220(.a(buffered_input), .b(12'b100010101100), .eq(weq2220));
    equaln #(12) e2221(.a(buffered_input), .b(12'b100010101101), .eq(weq2221));
    equaln #(12) e2222(.a(buffered_input), .b(12'b100010101110), .eq(weq2222));
    equaln #(12) e2223(.a(buffered_input), .b(12'b100010101111), .eq(weq2223));
    equaln #(12) e2224(.a(buffered_input), .b(12'b100010110000), .eq(weq2224));
    equaln #(12) e2225(.a(buffered_input), .b(12'b100010110001), .eq(weq2225));
    equaln #(12) e2226(.a(buffered_input), .b(12'b100010110010), .eq(weq2226));
    equaln #(12) e2227(.a(buffered_input), .b(12'b100010110011), .eq(weq2227));
    equaln #(12) e2228(.a(buffered_input), .b(12'b100010110100), .eq(weq2228));
    equaln #(12) e2229(.a(buffered_input), .b(12'b100010110101), .eq(weq2229));
    equaln #(12) e2230(.a(buffered_input), .b(12'b100010110110), .eq(weq2230));
    equaln #(12) e2231(.a(buffered_input), .b(12'b100010110111), .eq(weq2231));
    equaln #(12) e2232(.a(buffered_input), .b(12'b100010111000), .eq(weq2232));
    equaln #(12) e2233(.a(buffered_input), .b(12'b100010111001), .eq(weq2233));
    equaln #(12) e2234(.a(buffered_input), .b(12'b100010111010), .eq(weq2234));
    equaln #(12) e2235(.a(buffered_input), .b(12'b100010111011), .eq(weq2235));
    equaln #(12) e2236(.a(buffered_input), .b(12'b100010111100), .eq(weq2236));
    equaln #(12) e2237(.a(buffered_input), .b(12'b100010111101), .eq(weq2237));
    equaln #(12) e2238(.a(buffered_input), .b(12'b100010111110), .eq(weq2238));
    equaln #(12) e2239(.a(buffered_input), .b(12'b100010111111), .eq(weq2239));
    equaln #(12) e2240(.a(buffered_input), .b(12'b100011000000), .eq(weq2240));
    equaln #(12) e2241(.a(buffered_input), .b(12'b100011000001), .eq(weq2241));
    equaln #(12) e2242(.a(buffered_input), .b(12'b100011000010), .eq(weq2242));
    equaln #(12) e2243(.a(buffered_input), .b(12'b100011000011), .eq(weq2243));
    equaln #(12) e2244(.a(buffered_input), .b(12'b100011000100), .eq(weq2244));
    equaln #(12) e2245(.a(buffered_input), .b(12'b100011000101), .eq(weq2245));
    equaln #(12) e2246(.a(buffered_input), .b(12'b100011000110), .eq(weq2246));
    equaln #(12) e2247(.a(buffered_input), .b(12'b100011000111), .eq(weq2247));
    equaln #(12) e2248(.a(buffered_input), .b(12'b100011001000), .eq(weq2248));
    equaln #(12) e2249(.a(buffered_input), .b(12'b100011001001), .eq(weq2249));
    equaln #(12) e2250(.a(buffered_input), .b(12'b100011001010), .eq(weq2250));
    equaln #(12) e2251(.a(buffered_input), .b(12'b100011001011), .eq(weq2251));
    equaln #(12) e2252(.a(buffered_input), .b(12'b100011001100), .eq(weq2252));
    equaln #(12) e2253(.a(buffered_input), .b(12'b100011001101), .eq(weq2253));
    equaln #(12) e2254(.a(buffered_input), .b(12'b100011001110), .eq(weq2254));
    equaln #(12) e2255(.a(buffered_input), .b(12'b100011001111), .eq(weq2255));
    equaln #(12) e2256(.a(buffered_input), .b(12'b100011010000), .eq(weq2256));
    equaln #(12) e2257(.a(buffered_input), .b(12'b100011010001), .eq(weq2257));
    equaln #(12) e2258(.a(buffered_input), .b(12'b100011010010), .eq(weq2258));
    equaln #(12) e2259(.a(buffered_input), .b(12'b100011010011), .eq(weq2259));
    equaln #(12) e2260(.a(buffered_input), .b(12'b100011010100), .eq(weq2260));
    equaln #(12) e2261(.a(buffered_input), .b(12'b100011010101), .eq(weq2261));
    equaln #(12) e2262(.a(buffered_input), .b(12'b100011010110), .eq(weq2262));
    equaln #(12) e2263(.a(buffered_input), .b(12'b100011010111), .eq(weq2263));
    equaln #(12) e2264(.a(buffered_input), .b(12'b100011011000), .eq(weq2264));
    equaln #(12) e2265(.a(buffered_input), .b(12'b100011011001), .eq(weq2265));
    equaln #(12) e2266(.a(buffered_input), .b(12'b100011011010), .eq(weq2266));
    equaln #(12) e2267(.a(buffered_input), .b(12'b100011011011), .eq(weq2267));
    equaln #(12) e2268(.a(buffered_input), .b(12'b100011011100), .eq(weq2268));
    equaln #(12) e2269(.a(buffered_input), .b(12'b100011011101), .eq(weq2269));
    equaln #(12) e2270(.a(buffered_input), .b(12'b100011011110), .eq(weq2270));
    equaln #(12) e2271(.a(buffered_input), .b(12'b100011011111), .eq(weq2271));
    equaln #(12) e2272(.a(buffered_input), .b(12'b100011100000), .eq(weq2272));
    equaln #(12) e2273(.a(buffered_input), .b(12'b100011100001), .eq(weq2273));
    equaln #(12) e2274(.a(buffered_input), .b(12'b100011100010), .eq(weq2274));
    equaln #(12) e2275(.a(buffered_input), .b(12'b100011100011), .eq(weq2275));
    equaln #(12) e2276(.a(buffered_input), .b(12'b100011100100), .eq(weq2276));
    equaln #(12) e2277(.a(buffered_input), .b(12'b100011100101), .eq(weq2277));
    equaln #(12) e2278(.a(buffered_input), .b(12'b100011100110), .eq(weq2278));
    equaln #(12) e2279(.a(buffered_input), .b(12'b100011100111), .eq(weq2279));
    equaln #(12) e2280(.a(buffered_input), .b(12'b100011101000), .eq(weq2280));
    equaln #(12) e2281(.a(buffered_input), .b(12'b100011101001), .eq(weq2281));
    equaln #(12) e2282(.a(buffered_input), .b(12'b100011101010), .eq(weq2282));
    equaln #(12) e2283(.a(buffered_input), .b(12'b100011101011), .eq(weq2283));
    equaln #(12) e2284(.a(buffered_input), .b(12'b100011101100), .eq(weq2284));
    equaln #(12) e2285(.a(buffered_input), .b(12'b100011101101), .eq(weq2285));
    equaln #(12) e2286(.a(buffered_input), .b(12'b100011101110), .eq(weq2286));
    equaln #(12) e2287(.a(buffered_input), .b(12'b100011101111), .eq(weq2287));
    equaln #(12) e2288(.a(buffered_input), .b(12'b100011110000), .eq(weq2288));
    equaln #(12) e2289(.a(buffered_input), .b(12'b100011110001), .eq(weq2289));
    equaln #(12) e2290(.a(buffered_input), .b(12'b100011110010), .eq(weq2290));
    equaln #(12) e2291(.a(buffered_input), .b(12'b100011110011), .eq(weq2291));
    equaln #(12) e2292(.a(buffered_input), .b(12'b100011110100), .eq(weq2292));
    equaln #(12) e2293(.a(buffered_input), .b(12'b100011110101), .eq(weq2293));
    equaln #(12) e2294(.a(buffered_input), .b(12'b100011110110), .eq(weq2294));
    equaln #(12) e2295(.a(buffered_input), .b(12'b100011110111), .eq(weq2295));
    equaln #(12) e2296(.a(buffered_input), .b(12'b100011111000), .eq(weq2296));
    equaln #(12) e2297(.a(buffered_input), .b(12'b100011111001), .eq(weq2297));
    equaln #(12) e2298(.a(buffered_input), .b(12'b100011111010), .eq(weq2298));
    equaln #(12) e2299(.a(buffered_input), .b(12'b100011111011), .eq(weq2299));
    equaln #(12) e2300(.a(buffered_input), .b(12'b100011111100), .eq(weq2300));
    equaln #(12) e2301(.a(buffered_input), .b(12'b100011111101), .eq(weq2301));
    equaln #(12) e2302(.a(buffered_input), .b(12'b100011111110), .eq(weq2302));
    equaln #(12) e2303(.a(buffered_input), .b(12'b100011111111), .eq(weq2303));
    equaln #(12) e2304(.a(buffered_input), .b(12'b100100000000), .eq(weq2304));
    equaln #(12) e2305(.a(buffered_input), .b(12'b100100000001), .eq(weq2305));
    equaln #(12) e2306(.a(buffered_input), .b(12'b100100000010), .eq(weq2306));
    equaln #(12) e2307(.a(buffered_input), .b(12'b100100000011), .eq(weq2307));
    equaln #(12) e2308(.a(buffered_input), .b(12'b100100000100), .eq(weq2308));
    equaln #(12) e2309(.a(buffered_input), .b(12'b100100000101), .eq(weq2309));
    equaln #(12) e2310(.a(buffered_input), .b(12'b100100000110), .eq(weq2310));
    equaln #(12) e2311(.a(buffered_input), .b(12'b100100000111), .eq(weq2311));
    equaln #(12) e2312(.a(buffered_input), .b(12'b100100001000), .eq(weq2312));
    equaln #(12) e2313(.a(buffered_input), .b(12'b100100001001), .eq(weq2313));
    equaln #(12) e2314(.a(buffered_input), .b(12'b100100001010), .eq(weq2314));
    equaln #(12) e2315(.a(buffered_input), .b(12'b100100001011), .eq(weq2315));
    equaln #(12) e2316(.a(buffered_input), .b(12'b100100001100), .eq(weq2316));
    equaln #(12) e2317(.a(buffered_input), .b(12'b100100001101), .eq(weq2317));
    equaln #(12) e2318(.a(buffered_input), .b(12'b100100001110), .eq(weq2318));
    equaln #(12) e2319(.a(buffered_input), .b(12'b100100001111), .eq(weq2319));
    equaln #(12) e2320(.a(buffered_input), .b(12'b100100010000), .eq(weq2320));
    equaln #(12) e2321(.a(buffered_input), .b(12'b100100010001), .eq(weq2321));
    equaln #(12) e2322(.a(buffered_input), .b(12'b100100010010), .eq(weq2322));
    equaln #(12) e2323(.a(buffered_input), .b(12'b100100010011), .eq(weq2323));
    equaln #(12) e2324(.a(buffered_input), .b(12'b100100010100), .eq(weq2324));
    equaln #(12) e2325(.a(buffered_input), .b(12'b100100010101), .eq(weq2325));
    equaln #(12) e2326(.a(buffered_input), .b(12'b100100010110), .eq(weq2326));
    equaln #(12) e2327(.a(buffered_input), .b(12'b100100010111), .eq(weq2327));
    equaln #(12) e2328(.a(buffered_input), .b(12'b100100011000), .eq(weq2328));
    equaln #(12) e2329(.a(buffered_input), .b(12'b100100011001), .eq(weq2329));
    equaln #(12) e2330(.a(buffered_input), .b(12'b100100011010), .eq(weq2330));
    equaln #(12) e2331(.a(buffered_input), .b(12'b100100011011), .eq(weq2331));
    equaln #(12) e2332(.a(buffered_input), .b(12'b100100011100), .eq(weq2332));
    equaln #(12) e2333(.a(buffered_input), .b(12'b100100011101), .eq(weq2333));
    equaln #(12) e2334(.a(buffered_input), .b(12'b100100011110), .eq(weq2334));
    equaln #(12) e2335(.a(buffered_input), .b(12'b100100011111), .eq(weq2335));
    equaln #(12) e2336(.a(buffered_input), .b(12'b100100100000), .eq(weq2336));
    equaln #(12) e2337(.a(buffered_input), .b(12'b100100100001), .eq(weq2337));
    equaln #(12) e2338(.a(buffered_input), .b(12'b100100100010), .eq(weq2338));
    equaln #(12) e2339(.a(buffered_input), .b(12'b100100100011), .eq(weq2339));
    equaln #(12) e2340(.a(buffered_input), .b(12'b100100100100), .eq(weq2340));
    equaln #(12) e2341(.a(buffered_input), .b(12'b100100100101), .eq(weq2341));
    equaln #(12) e2342(.a(buffered_input), .b(12'b100100100110), .eq(weq2342));
    equaln #(12) e2343(.a(buffered_input), .b(12'b100100100111), .eq(weq2343));
    equaln #(12) e2344(.a(buffered_input), .b(12'b100100101000), .eq(weq2344));
    equaln #(12) e2345(.a(buffered_input), .b(12'b100100101001), .eq(weq2345));
    equaln #(12) e2346(.a(buffered_input), .b(12'b100100101010), .eq(weq2346));
    equaln #(12) e2347(.a(buffered_input), .b(12'b100100101011), .eq(weq2347));
    equaln #(12) e2348(.a(buffered_input), .b(12'b100100101100), .eq(weq2348));
    equaln #(12) e2349(.a(buffered_input), .b(12'b100100101101), .eq(weq2349));
    equaln #(12) e2350(.a(buffered_input), .b(12'b100100101110), .eq(weq2350));
    equaln #(12) e2351(.a(buffered_input), .b(12'b100100101111), .eq(weq2351));
    equaln #(12) e2352(.a(buffered_input), .b(12'b100100110000), .eq(weq2352));
    equaln #(12) e2353(.a(buffered_input), .b(12'b100100110001), .eq(weq2353));
    equaln #(12) e2354(.a(buffered_input), .b(12'b100100110010), .eq(weq2354));
    equaln #(12) e2355(.a(buffered_input), .b(12'b100100110011), .eq(weq2355));
    equaln #(12) e2356(.a(buffered_input), .b(12'b100100110100), .eq(weq2356));
    equaln #(12) e2357(.a(buffered_input), .b(12'b100100110101), .eq(weq2357));
    equaln #(12) e2358(.a(buffered_input), .b(12'b100100110110), .eq(weq2358));
    equaln #(12) e2359(.a(buffered_input), .b(12'b100100110111), .eq(weq2359));
    equaln #(12) e2360(.a(buffered_input), .b(12'b100100111000), .eq(weq2360));
    equaln #(12) e2361(.a(buffered_input), .b(12'b100100111001), .eq(weq2361));
    equaln #(12) e2362(.a(buffered_input), .b(12'b100100111010), .eq(weq2362));
    equaln #(12) e2363(.a(buffered_input), .b(12'b100100111011), .eq(weq2363));
    equaln #(12) e2364(.a(buffered_input), .b(12'b100100111100), .eq(weq2364));
    equaln #(12) e2365(.a(buffered_input), .b(12'b100100111101), .eq(weq2365));
    equaln #(12) e2366(.a(buffered_input), .b(12'b100100111110), .eq(weq2366));
    equaln #(12) e2367(.a(buffered_input), .b(12'b100100111111), .eq(weq2367));
    equaln #(12) e2368(.a(buffered_input), .b(12'b100101000000), .eq(weq2368));
    equaln #(12) e2369(.a(buffered_input), .b(12'b100101000001), .eq(weq2369));
    equaln #(12) e2370(.a(buffered_input), .b(12'b100101000010), .eq(weq2370));
    equaln #(12) e2371(.a(buffered_input), .b(12'b100101000011), .eq(weq2371));
    equaln #(12) e2372(.a(buffered_input), .b(12'b100101000100), .eq(weq2372));
    equaln #(12) e2373(.a(buffered_input), .b(12'b100101000101), .eq(weq2373));
    equaln #(12) e2374(.a(buffered_input), .b(12'b100101000110), .eq(weq2374));
    equaln #(12) e2375(.a(buffered_input), .b(12'b100101000111), .eq(weq2375));
    equaln #(12) e2376(.a(buffered_input), .b(12'b100101001000), .eq(weq2376));
    equaln #(12) e2377(.a(buffered_input), .b(12'b100101001001), .eq(weq2377));
    equaln #(12) e2378(.a(buffered_input), .b(12'b100101001010), .eq(weq2378));
    equaln #(12) e2379(.a(buffered_input), .b(12'b100101001011), .eq(weq2379));
    equaln #(12) e2380(.a(buffered_input), .b(12'b100101001100), .eq(weq2380));
    equaln #(12) e2381(.a(buffered_input), .b(12'b100101001101), .eq(weq2381));
    equaln #(12) e2382(.a(buffered_input), .b(12'b100101001110), .eq(weq2382));
    equaln #(12) e2383(.a(buffered_input), .b(12'b100101001111), .eq(weq2383));
    equaln #(12) e2384(.a(buffered_input), .b(12'b100101010000), .eq(weq2384));
    equaln #(12) e2385(.a(buffered_input), .b(12'b100101010001), .eq(weq2385));
    equaln #(12) e2386(.a(buffered_input), .b(12'b100101010010), .eq(weq2386));
    equaln #(12) e2387(.a(buffered_input), .b(12'b100101010011), .eq(weq2387));
    equaln #(12) e2388(.a(buffered_input), .b(12'b100101010100), .eq(weq2388));
    equaln #(12) e2389(.a(buffered_input), .b(12'b100101010101), .eq(weq2389));
    equaln #(12) e2390(.a(buffered_input), .b(12'b100101010110), .eq(weq2390));
    equaln #(12) e2391(.a(buffered_input), .b(12'b100101010111), .eq(weq2391));
    equaln #(12) e2392(.a(buffered_input), .b(12'b100101011000), .eq(weq2392));
    equaln #(12) e2393(.a(buffered_input), .b(12'b100101011001), .eq(weq2393));
    equaln #(12) e2394(.a(buffered_input), .b(12'b100101011010), .eq(weq2394));
    equaln #(12) e2395(.a(buffered_input), .b(12'b100101011011), .eq(weq2395));
    equaln #(12) e2396(.a(buffered_input), .b(12'b100101011100), .eq(weq2396));
    equaln #(12) e2397(.a(buffered_input), .b(12'b100101011101), .eq(weq2397));
    equaln #(12) e2398(.a(buffered_input), .b(12'b100101011110), .eq(weq2398));
    equaln #(12) e2399(.a(buffered_input), .b(12'b100101011111), .eq(weq2399));
    equaln #(12) e2400(.a(buffered_input), .b(12'b100101100000), .eq(weq2400));
    equaln #(12) e2401(.a(buffered_input), .b(12'b100101100001), .eq(weq2401));
    equaln #(12) e2402(.a(buffered_input), .b(12'b100101100010), .eq(weq2402));
    equaln #(12) e2403(.a(buffered_input), .b(12'b100101100011), .eq(weq2403));
    equaln #(12) e2404(.a(buffered_input), .b(12'b100101100100), .eq(weq2404));
    equaln #(12) e2405(.a(buffered_input), .b(12'b100101100101), .eq(weq2405));
    equaln #(12) e2406(.a(buffered_input), .b(12'b100101100110), .eq(weq2406));
    equaln #(12) e2407(.a(buffered_input), .b(12'b100101100111), .eq(weq2407));
    equaln #(12) e2408(.a(buffered_input), .b(12'b100101101000), .eq(weq2408));
    equaln #(12) e2409(.a(buffered_input), .b(12'b100101101001), .eq(weq2409));
    equaln #(12) e2410(.a(buffered_input), .b(12'b100101101010), .eq(weq2410));
    equaln #(12) e2411(.a(buffered_input), .b(12'b100101101011), .eq(weq2411));
    equaln #(12) e2412(.a(buffered_input), .b(12'b100101101100), .eq(weq2412));
    equaln #(12) e2413(.a(buffered_input), .b(12'b100101101101), .eq(weq2413));
    equaln #(12) e2414(.a(buffered_input), .b(12'b100101101110), .eq(weq2414));
    equaln #(12) e2415(.a(buffered_input), .b(12'b100101101111), .eq(weq2415));
    equaln #(12) e2416(.a(buffered_input), .b(12'b100101110000), .eq(weq2416));
    equaln #(12) e2417(.a(buffered_input), .b(12'b100101110001), .eq(weq2417));
    equaln #(12) e2418(.a(buffered_input), .b(12'b100101110010), .eq(weq2418));
    equaln #(12) e2419(.a(buffered_input), .b(12'b100101110011), .eq(weq2419));
    equaln #(12) e2420(.a(buffered_input), .b(12'b100101110100), .eq(weq2420));
    equaln #(12) e2421(.a(buffered_input), .b(12'b100101110101), .eq(weq2421));
    equaln #(12) e2422(.a(buffered_input), .b(12'b100101110110), .eq(weq2422));
    equaln #(12) e2423(.a(buffered_input), .b(12'b100101110111), .eq(weq2423));
    equaln #(12) e2424(.a(buffered_input), .b(12'b100101111000), .eq(weq2424));
    equaln #(12) e2425(.a(buffered_input), .b(12'b100101111001), .eq(weq2425));
    equaln #(12) e2426(.a(buffered_input), .b(12'b100101111010), .eq(weq2426));
    equaln #(12) e2427(.a(buffered_input), .b(12'b100101111011), .eq(weq2427));
    equaln #(12) e2428(.a(buffered_input), .b(12'b100101111100), .eq(weq2428));
    equaln #(12) e2429(.a(buffered_input), .b(12'b100101111101), .eq(weq2429));
    equaln #(12) e2430(.a(buffered_input), .b(12'b100101111110), .eq(weq2430));
    equaln #(12) e2431(.a(buffered_input), .b(12'b100101111111), .eq(weq2431));
    equaln #(12) e2432(.a(buffered_input), .b(12'b100110000000), .eq(weq2432));
    equaln #(12) e2433(.a(buffered_input), .b(12'b100110000001), .eq(weq2433));
    equaln #(12) e2434(.a(buffered_input), .b(12'b100110000010), .eq(weq2434));
    equaln #(12) e2435(.a(buffered_input), .b(12'b100110000011), .eq(weq2435));
    equaln #(12) e2436(.a(buffered_input), .b(12'b100110000100), .eq(weq2436));
    equaln #(12) e2437(.a(buffered_input), .b(12'b100110000101), .eq(weq2437));
    equaln #(12) e2438(.a(buffered_input), .b(12'b100110000110), .eq(weq2438));
    equaln #(12) e2439(.a(buffered_input), .b(12'b100110000111), .eq(weq2439));
    equaln #(12) e2440(.a(buffered_input), .b(12'b100110001000), .eq(weq2440));
    equaln #(12) e2441(.a(buffered_input), .b(12'b100110001001), .eq(weq2441));
    equaln #(12) e2442(.a(buffered_input), .b(12'b100110001010), .eq(weq2442));
    equaln #(12) e2443(.a(buffered_input), .b(12'b100110001011), .eq(weq2443));
    equaln #(12) e2444(.a(buffered_input), .b(12'b100110001100), .eq(weq2444));
    equaln #(12) e2445(.a(buffered_input), .b(12'b100110001101), .eq(weq2445));
    equaln #(12) e2446(.a(buffered_input), .b(12'b100110001110), .eq(weq2446));
    equaln #(12) e2447(.a(buffered_input), .b(12'b100110001111), .eq(weq2447));
    equaln #(12) e2448(.a(buffered_input), .b(12'b100110010000), .eq(weq2448));
    equaln #(12) e2449(.a(buffered_input), .b(12'b100110010001), .eq(weq2449));
    equaln #(12) e2450(.a(buffered_input), .b(12'b100110010010), .eq(weq2450));
    equaln #(12) e2451(.a(buffered_input), .b(12'b100110010011), .eq(weq2451));
    equaln #(12) e2452(.a(buffered_input), .b(12'b100110010100), .eq(weq2452));
    equaln #(12) e2453(.a(buffered_input), .b(12'b100110010101), .eq(weq2453));
    equaln #(12) e2454(.a(buffered_input), .b(12'b100110010110), .eq(weq2454));
    equaln #(12) e2455(.a(buffered_input), .b(12'b100110010111), .eq(weq2455));
    equaln #(12) e2456(.a(buffered_input), .b(12'b100110011000), .eq(weq2456));
    equaln #(12) e2457(.a(buffered_input), .b(12'b100110011001), .eq(weq2457));
    equaln #(12) e2458(.a(buffered_input), .b(12'b100110011010), .eq(weq2458));
    equaln #(12) e2459(.a(buffered_input), .b(12'b100110011011), .eq(weq2459));
    equaln #(12) e2460(.a(buffered_input), .b(12'b100110011100), .eq(weq2460));
    equaln #(12) e2461(.a(buffered_input), .b(12'b100110011101), .eq(weq2461));
    equaln #(12) e2462(.a(buffered_input), .b(12'b100110011110), .eq(weq2462));
    equaln #(12) e2463(.a(buffered_input), .b(12'b100110011111), .eq(weq2463));
    equaln #(12) e2464(.a(buffered_input), .b(12'b100110100000), .eq(weq2464));
    equaln #(12) e2465(.a(buffered_input), .b(12'b100110100001), .eq(weq2465));
    equaln #(12) e2466(.a(buffered_input), .b(12'b100110100010), .eq(weq2466));
    equaln #(12) e2467(.a(buffered_input), .b(12'b100110100011), .eq(weq2467));
    equaln #(12) e2468(.a(buffered_input), .b(12'b100110100100), .eq(weq2468));
    equaln #(12) e2469(.a(buffered_input), .b(12'b100110100101), .eq(weq2469));
    equaln #(12) e2470(.a(buffered_input), .b(12'b100110100110), .eq(weq2470));
    equaln #(12) e2471(.a(buffered_input), .b(12'b100110100111), .eq(weq2471));
    equaln #(12) e2472(.a(buffered_input), .b(12'b100110101000), .eq(weq2472));
    equaln #(12) e2473(.a(buffered_input), .b(12'b100110101001), .eq(weq2473));
    equaln #(12) e2474(.a(buffered_input), .b(12'b100110101010), .eq(weq2474));
    equaln #(12) e2475(.a(buffered_input), .b(12'b100110101011), .eq(weq2475));
    equaln #(12) e2476(.a(buffered_input), .b(12'b100110101100), .eq(weq2476));
    equaln #(12) e2477(.a(buffered_input), .b(12'b100110101101), .eq(weq2477));
    equaln #(12) e2478(.a(buffered_input), .b(12'b100110101110), .eq(weq2478));
    equaln #(12) e2479(.a(buffered_input), .b(12'b100110101111), .eq(weq2479));
    equaln #(12) e2480(.a(buffered_input), .b(12'b100110110000), .eq(weq2480));
    equaln #(12) e2481(.a(buffered_input), .b(12'b100110110001), .eq(weq2481));
    equaln #(12) e2482(.a(buffered_input), .b(12'b100110110010), .eq(weq2482));
    equaln #(12) e2483(.a(buffered_input), .b(12'b100110110011), .eq(weq2483));
    equaln #(12) e2484(.a(buffered_input), .b(12'b100110110100), .eq(weq2484));
    equaln #(12) e2485(.a(buffered_input), .b(12'b100110110101), .eq(weq2485));
    equaln #(12) e2486(.a(buffered_input), .b(12'b100110110110), .eq(weq2486));
    equaln #(12) e2487(.a(buffered_input), .b(12'b100110110111), .eq(weq2487));
    equaln #(12) e2488(.a(buffered_input), .b(12'b100110111000), .eq(weq2488));
    equaln #(12) e2489(.a(buffered_input), .b(12'b100110111001), .eq(weq2489));
    equaln #(12) e2490(.a(buffered_input), .b(12'b100110111010), .eq(weq2490));
    equaln #(12) e2491(.a(buffered_input), .b(12'b100110111011), .eq(weq2491));
    equaln #(12) e2492(.a(buffered_input), .b(12'b100110111100), .eq(weq2492));
    equaln #(12) e2493(.a(buffered_input), .b(12'b100110111101), .eq(weq2493));
    equaln #(12) e2494(.a(buffered_input), .b(12'b100110111110), .eq(weq2494));
    equaln #(12) e2495(.a(buffered_input), .b(12'b100110111111), .eq(weq2495));
    equaln #(12) e2496(.a(buffered_input), .b(12'b100111000000), .eq(weq2496));
    equaln #(12) e2497(.a(buffered_input), .b(12'b100111000001), .eq(weq2497));
    equaln #(12) e2498(.a(buffered_input), .b(12'b100111000010), .eq(weq2498));
    equaln #(12) e2499(.a(buffered_input), .b(12'b100111000011), .eq(weq2499));
    equaln #(12) e2500(.a(buffered_input), .b(12'b100111000100), .eq(weq2500));
    equaln #(12) e2501(.a(buffered_input), .b(12'b100111000101), .eq(weq2501));
    equaln #(12) e2502(.a(buffered_input), .b(12'b100111000110), .eq(weq2502));
    equaln #(12) e2503(.a(buffered_input), .b(12'b100111000111), .eq(weq2503));
    equaln #(12) e2504(.a(buffered_input), .b(12'b100111001000), .eq(weq2504));
    equaln #(12) e2505(.a(buffered_input), .b(12'b100111001001), .eq(weq2505));
    equaln #(12) e2506(.a(buffered_input), .b(12'b100111001010), .eq(weq2506));
    equaln #(12) e2507(.a(buffered_input), .b(12'b100111001011), .eq(weq2507));
    equaln #(12) e2508(.a(buffered_input), .b(12'b100111001100), .eq(weq2508));
    equaln #(12) e2509(.a(buffered_input), .b(12'b100111001101), .eq(weq2509));
    equaln #(12) e2510(.a(buffered_input), .b(12'b100111001110), .eq(weq2510));
    equaln #(12) e2511(.a(buffered_input), .b(12'b100111001111), .eq(weq2511));
    equaln #(12) e2512(.a(buffered_input), .b(12'b100111010000), .eq(weq2512));
    equaln #(12) e2513(.a(buffered_input), .b(12'b100111010001), .eq(weq2513));
    equaln #(12) e2514(.a(buffered_input), .b(12'b100111010010), .eq(weq2514));
    equaln #(12) e2515(.a(buffered_input), .b(12'b100111010011), .eq(weq2515));
    equaln #(12) e2516(.a(buffered_input), .b(12'b100111010100), .eq(weq2516));
    equaln #(12) e2517(.a(buffered_input), .b(12'b100111010101), .eq(weq2517));
    equaln #(12) e2518(.a(buffered_input), .b(12'b100111010110), .eq(weq2518));
    equaln #(12) e2519(.a(buffered_input), .b(12'b100111010111), .eq(weq2519));
    equaln #(12) e2520(.a(buffered_input), .b(12'b100111011000), .eq(weq2520));
    equaln #(12) e2521(.a(buffered_input), .b(12'b100111011001), .eq(weq2521));
    equaln #(12) e2522(.a(buffered_input), .b(12'b100111011010), .eq(weq2522));
    equaln #(12) e2523(.a(buffered_input), .b(12'b100111011011), .eq(weq2523));
    equaln #(12) e2524(.a(buffered_input), .b(12'b100111011100), .eq(weq2524));
    equaln #(12) e2525(.a(buffered_input), .b(12'b100111011101), .eq(weq2525));
    equaln #(12) e2526(.a(buffered_input), .b(12'b100111011110), .eq(weq2526));
    equaln #(12) e2527(.a(buffered_input), .b(12'b100111011111), .eq(weq2527));
    equaln #(12) e2528(.a(buffered_input), .b(12'b100111100000), .eq(weq2528));
    equaln #(12) e2529(.a(buffered_input), .b(12'b100111100001), .eq(weq2529));
    equaln #(12) e2530(.a(buffered_input), .b(12'b100111100010), .eq(weq2530));
    equaln #(12) e2531(.a(buffered_input), .b(12'b100111100011), .eq(weq2531));
    equaln #(12) e2532(.a(buffered_input), .b(12'b100111100100), .eq(weq2532));
    equaln #(12) e2533(.a(buffered_input), .b(12'b100111100101), .eq(weq2533));
    equaln #(12) e2534(.a(buffered_input), .b(12'b100111100110), .eq(weq2534));
    equaln #(12) e2535(.a(buffered_input), .b(12'b100111100111), .eq(weq2535));
    equaln #(12) e2536(.a(buffered_input), .b(12'b100111101000), .eq(weq2536));
    equaln #(12) e2537(.a(buffered_input), .b(12'b100111101001), .eq(weq2537));
    equaln #(12) e2538(.a(buffered_input), .b(12'b100111101010), .eq(weq2538));
    equaln #(12) e2539(.a(buffered_input), .b(12'b100111101011), .eq(weq2539));
    equaln #(12) e2540(.a(buffered_input), .b(12'b100111101100), .eq(weq2540));
    equaln #(12) e2541(.a(buffered_input), .b(12'b100111101101), .eq(weq2541));
    equaln #(12) e2542(.a(buffered_input), .b(12'b100111101110), .eq(weq2542));
    equaln #(12) e2543(.a(buffered_input), .b(12'b100111101111), .eq(weq2543));
    equaln #(12) e2544(.a(buffered_input), .b(12'b100111110000), .eq(weq2544));
    equaln #(12) e2545(.a(buffered_input), .b(12'b100111110001), .eq(weq2545));
    equaln #(12) e2546(.a(buffered_input), .b(12'b100111110010), .eq(weq2546));
    equaln #(12) e2547(.a(buffered_input), .b(12'b100111110011), .eq(weq2547));
    equaln #(12) e2548(.a(buffered_input), .b(12'b100111110100), .eq(weq2548));
    equaln #(12) e2549(.a(buffered_input), .b(12'b100111110101), .eq(weq2549));
    equaln #(12) e2550(.a(buffered_input), .b(12'b100111110110), .eq(weq2550));
    equaln #(12) e2551(.a(buffered_input), .b(12'b100111110111), .eq(weq2551));
    equaln #(12) e2552(.a(buffered_input), .b(12'b100111111000), .eq(weq2552));
    equaln #(12) e2553(.a(buffered_input), .b(12'b100111111001), .eq(weq2553));
    equaln #(12) e2554(.a(buffered_input), .b(12'b100111111010), .eq(weq2554));
    equaln #(12) e2555(.a(buffered_input), .b(12'b100111111011), .eq(weq2555));
    equaln #(12) e2556(.a(buffered_input), .b(12'b100111111100), .eq(weq2556));
    equaln #(12) e2557(.a(buffered_input), .b(12'b100111111101), .eq(weq2557));
    equaln #(12) e2558(.a(buffered_input), .b(12'b100111111110), .eq(weq2558));
    equaln #(12) e2559(.a(buffered_input), .b(12'b100111111111), .eq(weq2559));
    equaln #(12) e2560(.a(buffered_input), .b(12'b101000000000), .eq(weq2560));
    equaln #(12) e2561(.a(buffered_input), .b(12'b101000000001), .eq(weq2561));
    equaln #(12) e2562(.a(buffered_input), .b(12'b101000000010), .eq(weq2562));
    equaln #(12) e2563(.a(buffered_input), .b(12'b101000000011), .eq(weq2563));
    equaln #(12) e2564(.a(buffered_input), .b(12'b101000000100), .eq(weq2564));
    equaln #(12) e2565(.a(buffered_input), .b(12'b101000000101), .eq(weq2565));
    equaln #(12) e2566(.a(buffered_input), .b(12'b101000000110), .eq(weq2566));
    equaln #(12) e2567(.a(buffered_input), .b(12'b101000000111), .eq(weq2567));
    equaln #(12) e2568(.a(buffered_input), .b(12'b101000001000), .eq(weq2568));
    equaln #(12) e2569(.a(buffered_input), .b(12'b101000001001), .eq(weq2569));
    equaln #(12) e2570(.a(buffered_input), .b(12'b101000001010), .eq(weq2570));
    equaln #(12) e2571(.a(buffered_input), .b(12'b101000001011), .eq(weq2571));
    equaln #(12) e2572(.a(buffered_input), .b(12'b101000001100), .eq(weq2572));
    equaln #(12) e2573(.a(buffered_input), .b(12'b101000001101), .eq(weq2573));
    equaln #(12) e2574(.a(buffered_input), .b(12'b101000001110), .eq(weq2574));
    equaln #(12) e2575(.a(buffered_input), .b(12'b101000001111), .eq(weq2575));
    equaln #(12) e2576(.a(buffered_input), .b(12'b101000010000), .eq(weq2576));
    equaln #(12) e2577(.a(buffered_input), .b(12'b101000010001), .eq(weq2577));
    equaln #(12) e2578(.a(buffered_input), .b(12'b101000010010), .eq(weq2578));
    equaln #(12) e2579(.a(buffered_input), .b(12'b101000010011), .eq(weq2579));
    equaln #(12) e2580(.a(buffered_input), .b(12'b101000010100), .eq(weq2580));
    equaln #(12) e2581(.a(buffered_input), .b(12'b101000010101), .eq(weq2581));
    equaln #(12) e2582(.a(buffered_input), .b(12'b101000010110), .eq(weq2582));
    equaln #(12) e2583(.a(buffered_input), .b(12'b101000010111), .eq(weq2583));
    equaln #(12) e2584(.a(buffered_input), .b(12'b101000011000), .eq(weq2584));
    equaln #(12) e2585(.a(buffered_input), .b(12'b101000011001), .eq(weq2585));
    equaln #(12) e2586(.a(buffered_input), .b(12'b101000011010), .eq(weq2586));
    equaln #(12) e2587(.a(buffered_input), .b(12'b101000011011), .eq(weq2587));
    equaln #(12) e2588(.a(buffered_input), .b(12'b101000011100), .eq(weq2588));
    equaln #(12) e2589(.a(buffered_input), .b(12'b101000011101), .eq(weq2589));
    equaln #(12) e2590(.a(buffered_input), .b(12'b101000011110), .eq(weq2590));
    equaln #(12) e2591(.a(buffered_input), .b(12'b101000011111), .eq(weq2591));
    equaln #(12) e2592(.a(buffered_input), .b(12'b101000100000), .eq(weq2592));
    equaln #(12) e2593(.a(buffered_input), .b(12'b101000100001), .eq(weq2593));
    equaln #(12) e2594(.a(buffered_input), .b(12'b101000100010), .eq(weq2594));
    equaln #(12) e2595(.a(buffered_input), .b(12'b101000100011), .eq(weq2595));
    equaln #(12) e2596(.a(buffered_input), .b(12'b101000100100), .eq(weq2596));
    equaln #(12) e2597(.a(buffered_input), .b(12'b101000100101), .eq(weq2597));
    equaln #(12) e2598(.a(buffered_input), .b(12'b101000100110), .eq(weq2598));
    equaln #(12) e2599(.a(buffered_input), .b(12'b101000100111), .eq(weq2599));
    equaln #(12) e2600(.a(buffered_input), .b(12'b101000101000), .eq(weq2600));
    equaln #(12) e2601(.a(buffered_input), .b(12'b101000101001), .eq(weq2601));
    equaln #(12) e2602(.a(buffered_input), .b(12'b101000101010), .eq(weq2602));
    equaln #(12) e2603(.a(buffered_input), .b(12'b101000101011), .eq(weq2603));
    equaln #(12) e2604(.a(buffered_input), .b(12'b101000101100), .eq(weq2604));
    equaln #(12) e2605(.a(buffered_input), .b(12'b101000101101), .eq(weq2605));
    equaln #(12) e2606(.a(buffered_input), .b(12'b101000101110), .eq(weq2606));
    equaln #(12) e2607(.a(buffered_input), .b(12'b101000101111), .eq(weq2607));
    equaln #(12) e2608(.a(buffered_input), .b(12'b101000110000), .eq(weq2608));
    equaln #(12) e2609(.a(buffered_input), .b(12'b101000110001), .eq(weq2609));
    equaln #(12) e2610(.a(buffered_input), .b(12'b101000110010), .eq(weq2610));
    equaln #(12) e2611(.a(buffered_input), .b(12'b101000110011), .eq(weq2611));
    equaln #(12) e2612(.a(buffered_input), .b(12'b101000110100), .eq(weq2612));
    equaln #(12) e2613(.a(buffered_input), .b(12'b101000110101), .eq(weq2613));
    equaln #(12) e2614(.a(buffered_input), .b(12'b101000110110), .eq(weq2614));
    equaln #(12) e2615(.a(buffered_input), .b(12'b101000110111), .eq(weq2615));
    equaln #(12) e2616(.a(buffered_input), .b(12'b101000111000), .eq(weq2616));
    equaln #(12) e2617(.a(buffered_input), .b(12'b101000111001), .eq(weq2617));
    equaln #(12) e2618(.a(buffered_input), .b(12'b101000111010), .eq(weq2618));
    equaln #(12) e2619(.a(buffered_input), .b(12'b101000111011), .eq(weq2619));
    equaln #(12) e2620(.a(buffered_input), .b(12'b101000111100), .eq(weq2620));
    equaln #(12) e2621(.a(buffered_input), .b(12'b101000111101), .eq(weq2621));
    equaln #(12) e2622(.a(buffered_input), .b(12'b101000111110), .eq(weq2622));
    equaln #(12) e2623(.a(buffered_input), .b(12'b101000111111), .eq(weq2623));
    equaln #(12) e2624(.a(buffered_input), .b(12'b101001000000), .eq(weq2624));
    equaln #(12) e2625(.a(buffered_input), .b(12'b101001000001), .eq(weq2625));
    equaln #(12) e2626(.a(buffered_input), .b(12'b101001000010), .eq(weq2626));
    equaln #(12) e2627(.a(buffered_input), .b(12'b101001000011), .eq(weq2627));
    equaln #(12) e2628(.a(buffered_input), .b(12'b101001000100), .eq(weq2628));
    equaln #(12) e2629(.a(buffered_input), .b(12'b101001000101), .eq(weq2629));
    equaln #(12) e2630(.a(buffered_input), .b(12'b101001000110), .eq(weq2630));
    equaln #(12) e2631(.a(buffered_input), .b(12'b101001000111), .eq(weq2631));
    equaln #(12) e2632(.a(buffered_input), .b(12'b101001001000), .eq(weq2632));
    equaln #(12) e2633(.a(buffered_input), .b(12'b101001001001), .eq(weq2633));
    equaln #(12) e2634(.a(buffered_input), .b(12'b101001001010), .eq(weq2634));
    equaln #(12) e2635(.a(buffered_input), .b(12'b101001001011), .eq(weq2635));
    equaln #(12) e2636(.a(buffered_input), .b(12'b101001001100), .eq(weq2636));
    equaln #(12) e2637(.a(buffered_input), .b(12'b101001001101), .eq(weq2637));
    equaln #(12) e2638(.a(buffered_input), .b(12'b101001001110), .eq(weq2638));
    equaln #(12) e2639(.a(buffered_input), .b(12'b101001001111), .eq(weq2639));
    equaln #(12) e2640(.a(buffered_input), .b(12'b101001010000), .eq(weq2640));
    equaln #(12) e2641(.a(buffered_input), .b(12'b101001010001), .eq(weq2641));
    equaln #(12) e2642(.a(buffered_input), .b(12'b101001010010), .eq(weq2642));
    equaln #(12) e2643(.a(buffered_input), .b(12'b101001010011), .eq(weq2643));
    equaln #(12) e2644(.a(buffered_input), .b(12'b101001010100), .eq(weq2644));
    equaln #(12) e2645(.a(buffered_input), .b(12'b101001010101), .eq(weq2645));
    equaln #(12) e2646(.a(buffered_input), .b(12'b101001010110), .eq(weq2646));
    equaln #(12) e2647(.a(buffered_input), .b(12'b101001010111), .eq(weq2647));
    equaln #(12) e2648(.a(buffered_input), .b(12'b101001011000), .eq(weq2648));
    equaln #(12) e2649(.a(buffered_input), .b(12'b101001011001), .eq(weq2649));
    equaln #(12) e2650(.a(buffered_input), .b(12'b101001011010), .eq(weq2650));
    equaln #(12) e2651(.a(buffered_input), .b(12'b101001011011), .eq(weq2651));
    equaln #(12) e2652(.a(buffered_input), .b(12'b101001011100), .eq(weq2652));
    equaln #(12) e2653(.a(buffered_input), .b(12'b101001011101), .eq(weq2653));
    equaln #(12) e2654(.a(buffered_input), .b(12'b101001011110), .eq(weq2654));
    equaln #(12) e2655(.a(buffered_input), .b(12'b101001011111), .eq(weq2655));
    equaln #(12) e2656(.a(buffered_input), .b(12'b101001100000), .eq(weq2656));
    equaln #(12) e2657(.a(buffered_input), .b(12'b101001100001), .eq(weq2657));
    equaln #(12) e2658(.a(buffered_input), .b(12'b101001100010), .eq(weq2658));
    equaln #(12) e2659(.a(buffered_input), .b(12'b101001100011), .eq(weq2659));
    equaln #(12) e2660(.a(buffered_input), .b(12'b101001100100), .eq(weq2660));
    equaln #(12) e2661(.a(buffered_input), .b(12'b101001100101), .eq(weq2661));
    equaln #(12) e2662(.a(buffered_input), .b(12'b101001100110), .eq(weq2662));
    equaln #(12) e2663(.a(buffered_input), .b(12'b101001100111), .eq(weq2663));
    equaln #(12) e2664(.a(buffered_input), .b(12'b101001101000), .eq(weq2664));
    equaln #(12) e2665(.a(buffered_input), .b(12'b101001101001), .eq(weq2665));
    equaln #(12) e2666(.a(buffered_input), .b(12'b101001101010), .eq(weq2666));
    equaln #(12) e2667(.a(buffered_input), .b(12'b101001101011), .eq(weq2667));
    equaln #(12) e2668(.a(buffered_input), .b(12'b101001101100), .eq(weq2668));
    equaln #(12) e2669(.a(buffered_input), .b(12'b101001101101), .eq(weq2669));
    equaln #(12) e2670(.a(buffered_input), .b(12'b101001101110), .eq(weq2670));
    equaln #(12) e2671(.a(buffered_input), .b(12'b101001101111), .eq(weq2671));
    equaln #(12) e2672(.a(buffered_input), .b(12'b101001110000), .eq(weq2672));
    equaln #(12) e2673(.a(buffered_input), .b(12'b101001110001), .eq(weq2673));
    equaln #(12) e2674(.a(buffered_input), .b(12'b101001110010), .eq(weq2674));
    equaln #(12) e2675(.a(buffered_input), .b(12'b101001110011), .eq(weq2675));
    equaln #(12) e2676(.a(buffered_input), .b(12'b101001110100), .eq(weq2676));
    equaln #(12) e2677(.a(buffered_input), .b(12'b101001110101), .eq(weq2677));
    equaln #(12) e2678(.a(buffered_input), .b(12'b101001110110), .eq(weq2678));
    equaln #(12) e2679(.a(buffered_input), .b(12'b101001110111), .eq(weq2679));
    equaln #(12) e2680(.a(buffered_input), .b(12'b101001111000), .eq(weq2680));
    equaln #(12) e2681(.a(buffered_input), .b(12'b101001111001), .eq(weq2681));
    equaln #(12) e2682(.a(buffered_input), .b(12'b101001111010), .eq(weq2682));
    equaln #(12) e2683(.a(buffered_input), .b(12'b101001111011), .eq(weq2683));
    equaln #(12) e2684(.a(buffered_input), .b(12'b101001111100), .eq(weq2684));
    equaln #(12) e2685(.a(buffered_input), .b(12'b101001111101), .eq(weq2685));
    equaln #(12) e2686(.a(buffered_input), .b(12'b101001111110), .eq(weq2686));
    equaln #(12) e2687(.a(buffered_input), .b(12'b101001111111), .eq(weq2687));
    equaln #(12) e2688(.a(buffered_input), .b(12'b101010000000), .eq(weq2688));
    equaln #(12) e2689(.a(buffered_input), .b(12'b101010000001), .eq(weq2689));
    equaln #(12) e2690(.a(buffered_input), .b(12'b101010000010), .eq(weq2690));
    equaln #(12) e2691(.a(buffered_input), .b(12'b101010000011), .eq(weq2691));
    equaln #(12) e2692(.a(buffered_input), .b(12'b101010000100), .eq(weq2692));
    equaln #(12) e2693(.a(buffered_input), .b(12'b101010000101), .eq(weq2693));
    equaln #(12) e2694(.a(buffered_input), .b(12'b101010000110), .eq(weq2694));
    equaln #(12) e2695(.a(buffered_input), .b(12'b101010000111), .eq(weq2695));
    equaln #(12) e2696(.a(buffered_input), .b(12'b101010001000), .eq(weq2696));
    equaln #(12) e2697(.a(buffered_input), .b(12'b101010001001), .eq(weq2697));
    equaln #(12) e2698(.a(buffered_input), .b(12'b101010001010), .eq(weq2698));
    equaln #(12) e2699(.a(buffered_input), .b(12'b101010001011), .eq(weq2699));
    equaln #(12) e2700(.a(buffered_input), .b(12'b101010001100), .eq(weq2700));
    equaln #(12) e2701(.a(buffered_input), .b(12'b101010001101), .eq(weq2701));
    equaln #(12) e2702(.a(buffered_input), .b(12'b101010001110), .eq(weq2702));
    equaln #(12) e2703(.a(buffered_input), .b(12'b101010001111), .eq(weq2703));
    equaln #(12) e2704(.a(buffered_input), .b(12'b101010010000), .eq(weq2704));
    equaln #(12) e2705(.a(buffered_input), .b(12'b101010010001), .eq(weq2705));
    equaln #(12) e2706(.a(buffered_input), .b(12'b101010010010), .eq(weq2706));
    equaln #(12) e2707(.a(buffered_input), .b(12'b101010010011), .eq(weq2707));
    equaln #(12) e2708(.a(buffered_input), .b(12'b101010010100), .eq(weq2708));
    equaln #(12) e2709(.a(buffered_input), .b(12'b101010010101), .eq(weq2709));
    equaln #(12) e2710(.a(buffered_input), .b(12'b101010010110), .eq(weq2710));
    equaln #(12) e2711(.a(buffered_input), .b(12'b101010010111), .eq(weq2711));
    equaln #(12) e2712(.a(buffered_input), .b(12'b101010011000), .eq(weq2712));
    equaln #(12) e2713(.a(buffered_input), .b(12'b101010011001), .eq(weq2713));
    equaln #(12) e2714(.a(buffered_input), .b(12'b101010011010), .eq(weq2714));
    equaln #(12) e2715(.a(buffered_input), .b(12'b101010011011), .eq(weq2715));
    equaln #(12) e2716(.a(buffered_input), .b(12'b101010011100), .eq(weq2716));
    equaln #(12) e2717(.a(buffered_input), .b(12'b101010011101), .eq(weq2717));
    equaln #(12) e2718(.a(buffered_input), .b(12'b101010011110), .eq(weq2718));
    equaln #(12) e2719(.a(buffered_input), .b(12'b101010011111), .eq(weq2719));
    equaln #(12) e2720(.a(buffered_input), .b(12'b101010100000), .eq(weq2720));
    equaln #(12) e2721(.a(buffered_input), .b(12'b101010100001), .eq(weq2721));
    equaln #(12) e2722(.a(buffered_input), .b(12'b101010100010), .eq(weq2722));
    equaln #(12) e2723(.a(buffered_input), .b(12'b101010100011), .eq(weq2723));
    equaln #(12) e2724(.a(buffered_input), .b(12'b101010100100), .eq(weq2724));
    equaln #(12) e2725(.a(buffered_input), .b(12'b101010100101), .eq(weq2725));
    equaln #(12) e2726(.a(buffered_input), .b(12'b101010100110), .eq(weq2726));
    equaln #(12) e2727(.a(buffered_input), .b(12'b101010100111), .eq(weq2727));
    equaln #(12) e2728(.a(buffered_input), .b(12'b101010101000), .eq(weq2728));
    equaln #(12) e2729(.a(buffered_input), .b(12'b101010101001), .eq(weq2729));
    equaln #(12) e2730(.a(buffered_input), .b(12'b101010101010), .eq(weq2730));
    equaln #(12) e2731(.a(buffered_input), .b(12'b101010101011), .eq(weq2731));
    equaln #(12) e2732(.a(buffered_input), .b(12'b101010101100), .eq(weq2732));
    equaln #(12) e2733(.a(buffered_input), .b(12'b101010101101), .eq(weq2733));
    equaln #(12) e2734(.a(buffered_input), .b(12'b101010101110), .eq(weq2734));
    equaln #(12) e2735(.a(buffered_input), .b(12'b101010101111), .eq(weq2735));
    equaln #(12) e2736(.a(buffered_input), .b(12'b101010110000), .eq(weq2736));
    equaln #(12) e2737(.a(buffered_input), .b(12'b101010110001), .eq(weq2737));
    equaln #(12) e2738(.a(buffered_input), .b(12'b101010110010), .eq(weq2738));
    equaln #(12) e2739(.a(buffered_input), .b(12'b101010110011), .eq(weq2739));
    equaln #(12) e2740(.a(buffered_input), .b(12'b101010110100), .eq(weq2740));
    equaln #(12) e2741(.a(buffered_input), .b(12'b101010110101), .eq(weq2741));
    equaln #(12) e2742(.a(buffered_input), .b(12'b101010110110), .eq(weq2742));
    equaln #(12) e2743(.a(buffered_input), .b(12'b101010110111), .eq(weq2743));
    equaln #(12) e2744(.a(buffered_input), .b(12'b101010111000), .eq(weq2744));
    equaln #(12) e2745(.a(buffered_input), .b(12'b101010111001), .eq(weq2745));
    equaln #(12) e2746(.a(buffered_input), .b(12'b101010111010), .eq(weq2746));
    equaln #(12) e2747(.a(buffered_input), .b(12'b101010111011), .eq(weq2747));
    equaln #(12) e2748(.a(buffered_input), .b(12'b101010111100), .eq(weq2748));
    equaln #(12) e2749(.a(buffered_input), .b(12'b101010111101), .eq(weq2749));
    equaln #(12) e2750(.a(buffered_input), .b(12'b101010111110), .eq(weq2750));
    equaln #(12) e2751(.a(buffered_input), .b(12'b101010111111), .eq(weq2751));
    equaln #(12) e2752(.a(buffered_input), .b(12'b101011000000), .eq(weq2752));
    equaln #(12) e2753(.a(buffered_input), .b(12'b101011000001), .eq(weq2753));
    equaln #(12) e2754(.a(buffered_input), .b(12'b101011000010), .eq(weq2754));
    equaln #(12) e2755(.a(buffered_input), .b(12'b101011000011), .eq(weq2755));
    equaln #(12) e2756(.a(buffered_input), .b(12'b101011000100), .eq(weq2756));
    equaln #(12) e2757(.a(buffered_input), .b(12'b101011000101), .eq(weq2757));
    equaln #(12) e2758(.a(buffered_input), .b(12'b101011000110), .eq(weq2758));
    equaln #(12) e2759(.a(buffered_input), .b(12'b101011000111), .eq(weq2759));
    equaln #(12) e2760(.a(buffered_input), .b(12'b101011001000), .eq(weq2760));
    equaln #(12) e2761(.a(buffered_input), .b(12'b101011001001), .eq(weq2761));
    equaln #(12) e2762(.a(buffered_input), .b(12'b101011001010), .eq(weq2762));
    equaln #(12) e2763(.a(buffered_input), .b(12'b101011001011), .eq(weq2763));
    equaln #(12) e2764(.a(buffered_input), .b(12'b101011001100), .eq(weq2764));
    equaln #(12) e2765(.a(buffered_input), .b(12'b101011001101), .eq(weq2765));
    equaln #(12) e2766(.a(buffered_input), .b(12'b101011001110), .eq(weq2766));
    equaln #(12) e2767(.a(buffered_input), .b(12'b101011001111), .eq(weq2767));
    equaln #(12) e2768(.a(buffered_input), .b(12'b101011010000), .eq(weq2768));
    equaln #(12) e2769(.a(buffered_input), .b(12'b101011010001), .eq(weq2769));
    equaln #(12) e2770(.a(buffered_input), .b(12'b101011010010), .eq(weq2770));
    equaln #(12) e2771(.a(buffered_input), .b(12'b101011010011), .eq(weq2771));
    equaln #(12) e2772(.a(buffered_input), .b(12'b101011010100), .eq(weq2772));
    equaln #(12) e2773(.a(buffered_input), .b(12'b101011010101), .eq(weq2773));
    equaln #(12) e2774(.a(buffered_input), .b(12'b101011010110), .eq(weq2774));
    equaln #(12) e2775(.a(buffered_input), .b(12'b101011010111), .eq(weq2775));
    equaln #(12) e2776(.a(buffered_input), .b(12'b101011011000), .eq(weq2776));
    equaln #(12) e2777(.a(buffered_input), .b(12'b101011011001), .eq(weq2777));
    equaln #(12) e2778(.a(buffered_input), .b(12'b101011011010), .eq(weq2778));
    equaln #(12) e2779(.a(buffered_input), .b(12'b101011011011), .eq(weq2779));
    equaln #(12) e2780(.a(buffered_input), .b(12'b101011011100), .eq(weq2780));
    equaln #(12) e2781(.a(buffered_input), .b(12'b101011011101), .eq(weq2781));
    equaln #(12) e2782(.a(buffered_input), .b(12'b101011011110), .eq(weq2782));
    equaln #(12) e2783(.a(buffered_input), .b(12'b101011011111), .eq(weq2783));
    equaln #(12) e2784(.a(buffered_input), .b(12'b101011100000), .eq(weq2784));
    equaln #(12) e2785(.a(buffered_input), .b(12'b101011100001), .eq(weq2785));
    equaln #(12) e2786(.a(buffered_input), .b(12'b101011100010), .eq(weq2786));
    equaln #(12) e2787(.a(buffered_input), .b(12'b101011100011), .eq(weq2787));
    equaln #(12) e2788(.a(buffered_input), .b(12'b101011100100), .eq(weq2788));
    equaln #(12) e2789(.a(buffered_input), .b(12'b101011100101), .eq(weq2789));
    equaln #(12) e2790(.a(buffered_input), .b(12'b101011100110), .eq(weq2790));
    equaln #(12) e2791(.a(buffered_input), .b(12'b101011100111), .eq(weq2791));
    equaln #(12) e2792(.a(buffered_input), .b(12'b101011101000), .eq(weq2792));
    equaln #(12) e2793(.a(buffered_input), .b(12'b101011101001), .eq(weq2793));
    equaln #(12) e2794(.a(buffered_input), .b(12'b101011101010), .eq(weq2794));
    equaln #(12) e2795(.a(buffered_input), .b(12'b101011101011), .eq(weq2795));
    equaln #(12) e2796(.a(buffered_input), .b(12'b101011101100), .eq(weq2796));
    equaln #(12) e2797(.a(buffered_input), .b(12'b101011101101), .eq(weq2797));
    equaln #(12) e2798(.a(buffered_input), .b(12'b101011101110), .eq(weq2798));
    equaln #(12) e2799(.a(buffered_input), .b(12'b101011101111), .eq(weq2799));
    equaln #(12) e2800(.a(buffered_input), .b(12'b101011110000), .eq(weq2800));
    equaln #(12) e2801(.a(buffered_input), .b(12'b101011110001), .eq(weq2801));
    equaln #(12) e2802(.a(buffered_input), .b(12'b101011110010), .eq(weq2802));
    equaln #(12) e2803(.a(buffered_input), .b(12'b101011110011), .eq(weq2803));
    equaln #(12) e2804(.a(buffered_input), .b(12'b101011110100), .eq(weq2804));
    equaln #(12) e2805(.a(buffered_input), .b(12'b101011110101), .eq(weq2805));
    equaln #(12) e2806(.a(buffered_input), .b(12'b101011110110), .eq(weq2806));
    equaln #(12) e2807(.a(buffered_input), .b(12'b101011110111), .eq(weq2807));
    equaln #(12) e2808(.a(buffered_input), .b(12'b101011111000), .eq(weq2808));
    equaln #(12) e2809(.a(buffered_input), .b(12'b101011111001), .eq(weq2809));
    equaln #(12) e2810(.a(buffered_input), .b(12'b101011111010), .eq(weq2810));
    equaln #(12) e2811(.a(buffered_input), .b(12'b101011111011), .eq(weq2811));
    equaln #(12) e2812(.a(buffered_input), .b(12'b101011111100), .eq(weq2812));
    equaln #(12) e2813(.a(buffered_input), .b(12'b101011111101), .eq(weq2813));
    equaln #(12) e2814(.a(buffered_input), .b(12'b101011111110), .eq(weq2814));
    equaln #(12) e2815(.a(buffered_input), .b(12'b101011111111), .eq(weq2815));
    equaln #(12) e2816(.a(buffered_input), .b(12'b101100000000), .eq(weq2816));
    equaln #(12) e2817(.a(buffered_input), .b(12'b101100000001), .eq(weq2817));
    equaln #(12) e2818(.a(buffered_input), .b(12'b101100000010), .eq(weq2818));
    equaln #(12) e2819(.a(buffered_input), .b(12'b101100000011), .eq(weq2819));
    equaln #(12) e2820(.a(buffered_input), .b(12'b101100000100), .eq(weq2820));
    equaln #(12) e2821(.a(buffered_input), .b(12'b101100000101), .eq(weq2821));
    equaln #(12) e2822(.a(buffered_input), .b(12'b101100000110), .eq(weq2822));
    equaln #(12) e2823(.a(buffered_input), .b(12'b101100000111), .eq(weq2823));
    equaln #(12) e2824(.a(buffered_input), .b(12'b101100001000), .eq(weq2824));
    equaln #(12) e2825(.a(buffered_input), .b(12'b101100001001), .eq(weq2825));
    equaln #(12) e2826(.a(buffered_input), .b(12'b101100001010), .eq(weq2826));
    equaln #(12) e2827(.a(buffered_input), .b(12'b101100001011), .eq(weq2827));
    equaln #(12) e2828(.a(buffered_input), .b(12'b101100001100), .eq(weq2828));
    equaln #(12) e2829(.a(buffered_input), .b(12'b101100001101), .eq(weq2829));
    equaln #(12) e2830(.a(buffered_input), .b(12'b101100001110), .eq(weq2830));
    equaln #(12) e2831(.a(buffered_input), .b(12'b101100001111), .eq(weq2831));
    equaln #(12) e2832(.a(buffered_input), .b(12'b101100010000), .eq(weq2832));
    equaln #(12) e2833(.a(buffered_input), .b(12'b101100010001), .eq(weq2833));
    equaln #(12) e2834(.a(buffered_input), .b(12'b101100010010), .eq(weq2834));
    equaln #(12) e2835(.a(buffered_input), .b(12'b101100010011), .eq(weq2835));
    equaln #(12) e2836(.a(buffered_input), .b(12'b101100010100), .eq(weq2836));
    equaln #(12) e2837(.a(buffered_input), .b(12'b101100010101), .eq(weq2837));
    equaln #(12) e2838(.a(buffered_input), .b(12'b101100010110), .eq(weq2838));
    equaln #(12) e2839(.a(buffered_input), .b(12'b101100010111), .eq(weq2839));
    equaln #(12) e2840(.a(buffered_input), .b(12'b101100011000), .eq(weq2840));
    equaln #(12) e2841(.a(buffered_input), .b(12'b101100011001), .eq(weq2841));
    equaln #(12) e2842(.a(buffered_input), .b(12'b101100011010), .eq(weq2842));
    equaln #(12) e2843(.a(buffered_input), .b(12'b101100011011), .eq(weq2843));
    equaln #(12) e2844(.a(buffered_input), .b(12'b101100011100), .eq(weq2844));
    equaln #(12) e2845(.a(buffered_input), .b(12'b101100011101), .eq(weq2845));
    equaln #(12) e2846(.a(buffered_input), .b(12'b101100011110), .eq(weq2846));
    equaln #(12) e2847(.a(buffered_input), .b(12'b101100011111), .eq(weq2847));
    equaln #(12) e2848(.a(buffered_input), .b(12'b101100100000), .eq(weq2848));
    equaln #(12) e2849(.a(buffered_input), .b(12'b101100100001), .eq(weq2849));
    equaln #(12) e2850(.a(buffered_input), .b(12'b101100100010), .eq(weq2850));
    equaln #(12) e2851(.a(buffered_input), .b(12'b101100100011), .eq(weq2851));
    equaln #(12) e2852(.a(buffered_input), .b(12'b101100100100), .eq(weq2852));
    equaln #(12) e2853(.a(buffered_input), .b(12'b101100100101), .eq(weq2853));
    equaln #(12) e2854(.a(buffered_input), .b(12'b101100100110), .eq(weq2854));
    equaln #(12) e2855(.a(buffered_input), .b(12'b101100100111), .eq(weq2855));
    equaln #(12) e2856(.a(buffered_input), .b(12'b101100101000), .eq(weq2856));
    equaln #(12) e2857(.a(buffered_input), .b(12'b101100101001), .eq(weq2857));
    equaln #(12) e2858(.a(buffered_input), .b(12'b101100101010), .eq(weq2858));
    equaln #(12) e2859(.a(buffered_input), .b(12'b101100101011), .eq(weq2859));
    equaln #(12) e2860(.a(buffered_input), .b(12'b101100101100), .eq(weq2860));
    equaln #(12) e2861(.a(buffered_input), .b(12'b101100101101), .eq(weq2861));
    equaln #(12) e2862(.a(buffered_input), .b(12'b101100101110), .eq(weq2862));
    equaln #(12) e2863(.a(buffered_input), .b(12'b101100101111), .eq(weq2863));
    equaln #(12) e2864(.a(buffered_input), .b(12'b101100110000), .eq(weq2864));
    equaln #(12) e2865(.a(buffered_input), .b(12'b101100110001), .eq(weq2865));
    equaln #(12) e2866(.a(buffered_input), .b(12'b101100110010), .eq(weq2866));
    equaln #(12) e2867(.a(buffered_input), .b(12'b101100110011), .eq(weq2867));
    equaln #(12) e2868(.a(buffered_input), .b(12'b101100110100), .eq(weq2868));
    equaln #(12) e2869(.a(buffered_input), .b(12'b101100110101), .eq(weq2869));
    equaln #(12) e2870(.a(buffered_input), .b(12'b101100110110), .eq(weq2870));
    equaln #(12) e2871(.a(buffered_input), .b(12'b101100110111), .eq(weq2871));
    equaln #(12) e2872(.a(buffered_input), .b(12'b101100111000), .eq(weq2872));
    equaln #(12) e2873(.a(buffered_input), .b(12'b101100111001), .eq(weq2873));
    equaln #(12) e2874(.a(buffered_input), .b(12'b101100111010), .eq(weq2874));
    equaln #(12) e2875(.a(buffered_input), .b(12'b101100111011), .eq(weq2875));
    equaln #(12) e2876(.a(buffered_input), .b(12'b101100111100), .eq(weq2876));
    equaln #(12) e2877(.a(buffered_input), .b(12'b101100111101), .eq(weq2877));
    equaln #(12) e2878(.a(buffered_input), .b(12'b101100111110), .eq(weq2878));
    equaln #(12) e2879(.a(buffered_input), .b(12'b101100111111), .eq(weq2879));
    equaln #(12) e2880(.a(buffered_input), .b(12'b101101000000), .eq(weq2880));
    equaln #(12) e2881(.a(buffered_input), .b(12'b101101000001), .eq(weq2881));
    equaln #(12) e2882(.a(buffered_input), .b(12'b101101000010), .eq(weq2882));
    equaln #(12) e2883(.a(buffered_input), .b(12'b101101000011), .eq(weq2883));
    equaln #(12) e2884(.a(buffered_input), .b(12'b101101000100), .eq(weq2884));
    equaln #(12) e2885(.a(buffered_input), .b(12'b101101000101), .eq(weq2885));
    equaln #(12) e2886(.a(buffered_input), .b(12'b101101000110), .eq(weq2886));
    equaln #(12) e2887(.a(buffered_input), .b(12'b101101000111), .eq(weq2887));
    equaln #(12) e2888(.a(buffered_input), .b(12'b101101001000), .eq(weq2888));
    equaln #(12) e2889(.a(buffered_input), .b(12'b101101001001), .eq(weq2889));
    equaln #(12) e2890(.a(buffered_input), .b(12'b101101001010), .eq(weq2890));
    equaln #(12) e2891(.a(buffered_input), .b(12'b101101001011), .eq(weq2891));
    equaln #(12) e2892(.a(buffered_input), .b(12'b101101001100), .eq(weq2892));
    equaln #(12) e2893(.a(buffered_input), .b(12'b101101001101), .eq(weq2893));
    equaln #(12) e2894(.a(buffered_input), .b(12'b101101001110), .eq(weq2894));
    equaln #(12) e2895(.a(buffered_input), .b(12'b101101001111), .eq(weq2895));
    equaln #(12) e2896(.a(buffered_input), .b(12'b101101010000), .eq(weq2896));
    equaln #(12) e2897(.a(buffered_input), .b(12'b101101010001), .eq(weq2897));
    equaln #(12) e2898(.a(buffered_input), .b(12'b101101010010), .eq(weq2898));
    equaln #(12) e2899(.a(buffered_input), .b(12'b101101010011), .eq(weq2899));
    equaln #(12) e2900(.a(buffered_input), .b(12'b101101010100), .eq(weq2900));
    equaln #(12) e2901(.a(buffered_input), .b(12'b101101010101), .eq(weq2901));
    equaln #(12) e2902(.a(buffered_input), .b(12'b101101010110), .eq(weq2902));
    equaln #(12) e2903(.a(buffered_input), .b(12'b101101010111), .eq(weq2903));
    equaln #(12) e2904(.a(buffered_input), .b(12'b101101011000), .eq(weq2904));
    equaln #(12) e2905(.a(buffered_input), .b(12'b101101011001), .eq(weq2905));
    equaln #(12) e2906(.a(buffered_input), .b(12'b101101011010), .eq(weq2906));
    equaln #(12) e2907(.a(buffered_input), .b(12'b101101011011), .eq(weq2907));
    equaln #(12) e2908(.a(buffered_input), .b(12'b101101011100), .eq(weq2908));
    equaln #(12) e2909(.a(buffered_input), .b(12'b101101011101), .eq(weq2909));
    equaln #(12) e2910(.a(buffered_input), .b(12'b101101011110), .eq(weq2910));
    equaln #(12) e2911(.a(buffered_input), .b(12'b101101011111), .eq(weq2911));
    equaln #(12) e2912(.a(buffered_input), .b(12'b101101100000), .eq(weq2912));
    equaln #(12) e2913(.a(buffered_input), .b(12'b101101100001), .eq(weq2913));
    equaln #(12) e2914(.a(buffered_input), .b(12'b101101100010), .eq(weq2914));
    equaln #(12) e2915(.a(buffered_input), .b(12'b101101100011), .eq(weq2915));
    equaln #(12) e2916(.a(buffered_input), .b(12'b101101100100), .eq(weq2916));
    equaln #(12) e2917(.a(buffered_input), .b(12'b101101100101), .eq(weq2917));
    equaln #(12) e2918(.a(buffered_input), .b(12'b101101100110), .eq(weq2918));
    equaln #(12) e2919(.a(buffered_input), .b(12'b101101100111), .eq(weq2919));
    equaln #(12) e2920(.a(buffered_input), .b(12'b101101101000), .eq(weq2920));
    equaln #(12) e2921(.a(buffered_input), .b(12'b101101101001), .eq(weq2921));
    equaln #(12) e2922(.a(buffered_input), .b(12'b101101101010), .eq(weq2922));
    equaln #(12) e2923(.a(buffered_input), .b(12'b101101101011), .eq(weq2923));
    equaln #(12) e2924(.a(buffered_input), .b(12'b101101101100), .eq(weq2924));
    equaln #(12) e2925(.a(buffered_input), .b(12'b101101101101), .eq(weq2925));
    equaln #(12) e2926(.a(buffered_input), .b(12'b101101101110), .eq(weq2926));
    equaln #(12) e2927(.a(buffered_input), .b(12'b101101101111), .eq(weq2927));
    equaln #(12) e2928(.a(buffered_input), .b(12'b101101110000), .eq(weq2928));
    equaln #(12) e2929(.a(buffered_input), .b(12'b101101110001), .eq(weq2929));
    equaln #(12) e2930(.a(buffered_input), .b(12'b101101110010), .eq(weq2930));
    equaln #(12) e2931(.a(buffered_input), .b(12'b101101110011), .eq(weq2931));
    equaln #(12) e2932(.a(buffered_input), .b(12'b101101110100), .eq(weq2932));
    equaln #(12) e2933(.a(buffered_input), .b(12'b101101110101), .eq(weq2933));
    equaln #(12) e2934(.a(buffered_input), .b(12'b101101110110), .eq(weq2934));
    equaln #(12) e2935(.a(buffered_input), .b(12'b101101110111), .eq(weq2935));
    equaln #(12) e2936(.a(buffered_input), .b(12'b101101111000), .eq(weq2936));
    equaln #(12) e2937(.a(buffered_input), .b(12'b101101111001), .eq(weq2937));
    equaln #(12) e2938(.a(buffered_input), .b(12'b101101111010), .eq(weq2938));
    equaln #(12) e2939(.a(buffered_input), .b(12'b101101111011), .eq(weq2939));
    equaln #(12) e2940(.a(buffered_input), .b(12'b101101111100), .eq(weq2940));
    equaln #(12) e2941(.a(buffered_input), .b(12'b101101111101), .eq(weq2941));
    equaln #(12) e2942(.a(buffered_input), .b(12'b101101111110), .eq(weq2942));
    equaln #(12) e2943(.a(buffered_input), .b(12'b101101111111), .eq(weq2943));
    equaln #(12) e2944(.a(buffered_input), .b(12'b101110000000), .eq(weq2944));
    equaln #(12) e2945(.a(buffered_input), .b(12'b101110000001), .eq(weq2945));
    equaln #(12) e2946(.a(buffered_input), .b(12'b101110000010), .eq(weq2946));
    equaln #(12) e2947(.a(buffered_input), .b(12'b101110000011), .eq(weq2947));
    equaln #(12) e2948(.a(buffered_input), .b(12'b101110000100), .eq(weq2948));
    equaln #(12) e2949(.a(buffered_input), .b(12'b101110000101), .eq(weq2949));
    equaln #(12) e2950(.a(buffered_input), .b(12'b101110000110), .eq(weq2950));
    equaln #(12) e2951(.a(buffered_input), .b(12'b101110000111), .eq(weq2951));
    equaln #(12) e2952(.a(buffered_input), .b(12'b101110001000), .eq(weq2952));
    equaln #(12) e2953(.a(buffered_input), .b(12'b101110001001), .eq(weq2953));
    equaln #(12) e2954(.a(buffered_input), .b(12'b101110001010), .eq(weq2954));
    equaln #(12) e2955(.a(buffered_input), .b(12'b101110001011), .eq(weq2955));
    equaln #(12) e2956(.a(buffered_input), .b(12'b101110001100), .eq(weq2956));
    equaln #(12) e2957(.a(buffered_input), .b(12'b101110001101), .eq(weq2957));
    equaln #(12) e2958(.a(buffered_input), .b(12'b101110001110), .eq(weq2958));
    equaln #(12) e2959(.a(buffered_input), .b(12'b101110001111), .eq(weq2959));
    equaln #(12) e2960(.a(buffered_input), .b(12'b101110010000), .eq(weq2960));
    equaln #(12) e2961(.a(buffered_input), .b(12'b101110010001), .eq(weq2961));
    equaln #(12) e2962(.a(buffered_input), .b(12'b101110010010), .eq(weq2962));
    equaln #(12) e2963(.a(buffered_input), .b(12'b101110010011), .eq(weq2963));
    equaln #(12) e2964(.a(buffered_input), .b(12'b101110010100), .eq(weq2964));
    equaln #(12) e2965(.a(buffered_input), .b(12'b101110010101), .eq(weq2965));
    equaln #(12) e2966(.a(buffered_input), .b(12'b101110010110), .eq(weq2966));
    equaln #(12) e2967(.a(buffered_input), .b(12'b101110010111), .eq(weq2967));
    equaln #(12) e2968(.a(buffered_input), .b(12'b101110011000), .eq(weq2968));
    equaln #(12) e2969(.a(buffered_input), .b(12'b101110011001), .eq(weq2969));
    equaln #(12) e2970(.a(buffered_input), .b(12'b101110011010), .eq(weq2970));
    equaln #(12) e2971(.a(buffered_input), .b(12'b101110011011), .eq(weq2971));
    equaln #(12) e2972(.a(buffered_input), .b(12'b101110011100), .eq(weq2972));
    equaln #(12) e2973(.a(buffered_input), .b(12'b101110011101), .eq(weq2973));
    equaln #(12) e2974(.a(buffered_input), .b(12'b101110011110), .eq(weq2974));
    equaln #(12) e2975(.a(buffered_input), .b(12'b101110011111), .eq(weq2975));
    equaln #(12) e2976(.a(buffered_input), .b(12'b101110100000), .eq(weq2976));
    equaln #(12) e2977(.a(buffered_input), .b(12'b101110100001), .eq(weq2977));
    equaln #(12) e2978(.a(buffered_input), .b(12'b101110100010), .eq(weq2978));
    equaln #(12) e2979(.a(buffered_input), .b(12'b101110100011), .eq(weq2979));
    equaln #(12) e2980(.a(buffered_input), .b(12'b101110100100), .eq(weq2980));
    equaln #(12) e2981(.a(buffered_input), .b(12'b101110100101), .eq(weq2981));
    equaln #(12) e2982(.a(buffered_input), .b(12'b101110100110), .eq(weq2982));
    equaln #(12) e2983(.a(buffered_input), .b(12'b101110100111), .eq(weq2983));
    equaln #(12) e2984(.a(buffered_input), .b(12'b101110101000), .eq(weq2984));
    equaln #(12) e2985(.a(buffered_input), .b(12'b101110101001), .eq(weq2985));
    equaln #(12) e2986(.a(buffered_input), .b(12'b101110101010), .eq(weq2986));
    equaln #(12) e2987(.a(buffered_input), .b(12'b101110101011), .eq(weq2987));
    equaln #(12) e2988(.a(buffered_input), .b(12'b101110101100), .eq(weq2988));
    equaln #(12) e2989(.a(buffered_input), .b(12'b101110101101), .eq(weq2989));
    equaln #(12) e2990(.a(buffered_input), .b(12'b101110101110), .eq(weq2990));
    equaln #(12) e2991(.a(buffered_input), .b(12'b101110101111), .eq(weq2991));
    equaln #(12) e2992(.a(buffered_input), .b(12'b101110110000), .eq(weq2992));
    equaln #(12) e2993(.a(buffered_input), .b(12'b101110110001), .eq(weq2993));
    equaln #(12) e2994(.a(buffered_input), .b(12'b101110110010), .eq(weq2994));
    equaln #(12) e2995(.a(buffered_input), .b(12'b101110110011), .eq(weq2995));
    equaln #(12) e2996(.a(buffered_input), .b(12'b101110110100), .eq(weq2996));
    equaln #(12) e2997(.a(buffered_input), .b(12'b101110110101), .eq(weq2997));
    equaln #(12) e2998(.a(buffered_input), .b(12'b101110110110), .eq(weq2998));
    equaln #(12) e2999(.a(buffered_input), .b(12'b101110110111), .eq(weq2999));
    equaln #(12) e3000(.a(buffered_input), .b(12'b101110111000), .eq(weq3000));
    equaln #(12) e3001(.a(buffered_input), .b(12'b101110111001), .eq(weq3001));
    equaln #(12) e3002(.a(buffered_input), .b(12'b101110111010), .eq(weq3002));
    equaln #(12) e3003(.a(buffered_input), .b(12'b101110111011), .eq(weq3003));
    equaln #(12) e3004(.a(buffered_input), .b(12'b101110111100), .eq(weq3004));
    equaln #(12) e3005(.a(buffered_input), .b(12'b101110111101), .eq(weq3005));
    equaln #(12) e3006(.a(buffered_input), .b(12'b101110111110), .eq(weq3006));
    equaln #(12) e3007(.a(buffered_input), .b(12'b101110111111), .eq(weq3007));
    equaln #(12) e3008(.a(buffered_input), .b(12'b101111000000), .eq(weq3008));
    equaln #(12) e3009(.a(buffered_input), .b(12'b101111000001), .eq(weq3009));
    equaln #(12) e3010(.a(buffered_input), .b(12'b101111000010), .eq(weq3010));
    equaln #(12) e3011(.a(buffered_input), .b(12'b101111000011), .eq(weq3011));
    equaln #(12) e3012(.a(buffered_input), .b(12'b101111000100), .eq(weq3012));
    equaln #(12) e3013(.a(buffered_input), .b(12'b101111000101), .eq(weq3013));
    equaln #(12) e3014(.a(buffered_input), .b(12'b101111000110), .eq(weq3014));
    equaln #(12) e3015(.a(buffered_input), .b(12'b101111000111), .eq(weq3015));
    equaln #(12) e3016(.a(buffered_input), .b(12'b101111001000), .eq(weq3016));
    equaln #(12) e3017(.a(buffered_input), .b(12'b101111001001), .eq(weq3017));
    equaln #(12) e3018(.a(buffered_input), .b(12'b101111001010), .eq(weq3018));
    equaln #(12) e3019(.a(buffered_input), .b(12'b101111001011), .eq(weq3019));
    equaln #(12) e3020(.a(buffered_input), .b(12'b101111001100), .eq(weq3020));
    equaln #(12) e3021(.a(buffered_input), .b(12'b101111001101), .eq(weq3021));
    equaln #(12) e3022(.a(buffered_input), .b(12'b101111001110), .eq(weq3022));
    equaln #(12) e3023(.a(buffered_input), .b(12'b101111001111), .eq(weq3023));
    equaln #(12) e3024(.a(buffered_input), .b(12'b101111010000), .eq(weq3024));
    equaln #(12) e3025(.a(buffered_input), .b(12'b101111010001), .eq(weq3025));
    equaln #(12) e3026(.a(buffered_input), .b(12'b101111010010), .eq(weq3026));
    equaln #(12) e3027(.a(buffered_input), .b(12'b101111010011), .eq(weq3027));
    equaln #(12) e3028(.a(buffered_input), .b(12'b101111010100), .eq(weq3028));
    equaln #(12) e3029(.a(buffered_input), .b(12'b101111010101), .eq(weq3029));
    equaln #(12) e3030(.a(buffered_input), .b(12'b101111010110), .eq(weq3030));
    equaln #(12) e3031(.a(buffered_input), .b(12'b101111010111), .eq(weq3031));
    equaln #(12) e3032(.a(buffered_input), .b(12'b101111011000), .eq(weq3032));
    equaln #(12) e3033(.a(buffered_input), .b(12'b101111011001), .eq(weq3033));
    equaln #(12) e3034(.a(buffered_input), .b(12'b101111011010), .eq(weq3034));
    equaln #(12) e3035(.a(buffered_input), .b(12'b101111011011), .eq(weq3035));
    equaln #(12) e3036(.a(buffered_input), .b(12'b101111011100), .eq(weq3036));
    equaln #(12) e3037(.a(buffered_input), .b(12'b101111011101), .eq(weq3037));
    equaln #(12) e3038(.a(buffered_input), .b(12'b101111011110), .eq(weq3038));
    equaln #(12) e3039(.a(buffered_input), .b(12'b101111011111), .eq(weq3039));
    equaln #(12) e3040(.a(buffered_input), .b(12'b101111100000), .eq(weq3040));
    equaln #(12) e3041(.a(buffered_input), .b(12'b101111100001), .eq(weq3041));
    equaln #(12) e3042(.a(buffered_input), .b(12'b101111100010), .eq(weq3042));
    equaln #(12) e3043(.a(buffered_input), .b(12'b101111100011), .eq(weq3043));
    equaln #(12) e3044(.a(buffered_input), .b(12'b101111100100), .eq(weq3044));
    equaln #(12) e3045(.a(buffered_input), .b(12'b101111100101), .eq(weq3045));
    equaln #(12) e3046(.a(buffered_input), .b(12'b101111100110), .eq(weq3046));
    equaln #(12) e3047(.a(buffered_input), .b(12'b101111100111), .eq(weq3047));
    equaln #(12) e3048(.a(buffered_input), .b(12'b101111101000), .eq(weq3048));
    equaln #(12) e3049(.a(buffered_input), .b(12'b101111101001), .eq(weq3049));
    equaln #(12) e3050(.a(buffered_input), .b(12'b101111101010), .eq(weq3050));
    equaln #(12) e3051(.a(buffered_input), .b(12'b101111101011), .eq(weq3051));
    equaln #(12) e3052(.a(buffered_input), .b(12'b101111101100), .eq(weq3052));
    equaln #(12) e3053(.a(buffered_input), .b(12'b101111101101), .eq(weq3053));
    equaln #(12) e3054(.a(buffered_input), .b(12'b101111101110), .eq(weq3054));
    equaln #(12) e3055(.a(buffered_input), .b(12'b101111101111), .eq(weq3055));
    equaln #(12) e3056(.a(buffered_input), .b(12'b101111110000), .eq(weq3056));
    equaln #(12) e3057(.a(buffered_input), .b(12'b101111110001), .eq(weq3057));
    equaln #(12) e3058(.a(buffered_input), .b(12'b101111110010), .eq(weq3058));
    equaln #(12) e3059(.a(buffered_input), .b(12'b101111110011), .eq(weq3059));
    equaln #(12) e3060(.a(buffered_input), .b(12'b101111110100), .eq(weq3060));
    equaln #(12) e3061(.a(buffered_input), .b(12'b101111110101), .eq(weq3061));
    equaln #(12) e3062(.a(buffered_input), .b(12'b101111110110), .eq(weq3062));
    equaln #(12) e3063(.a(buffered_input), .b(12'b101111110111), .eq(weq3063));
    equaln #(12) e3064(.a(buffered_input), .b(12'b101111111000), .eq(weq3064));
    equaln #(12) e3065(.a(buffered_input), .b(12'b101111111001), .eq(weq3065));
    equaln #(12) e3066(.a(buffered_input), .b(12'b101111111010), .eq(weq3066));
    equaln #(12) e3067(.a(buffered_input), .b(12'b101111111011), .eq(weq3067));
    equaln #(12) e3068(.a(buffered_input), .b(12'b101111111100), .eq(weq3068));
    equaln #(12) e3069(.a(buffered_input), .b(12'b101111111101), .eq(weq3069));
    equaln #(12) e3070(.a(buffered_input), .b(12'b101111111110), .eq(weq3070));
    equaln #(12) e3071(.a(buffered_input), .b(12'b101111111111), .eq(weq3071));
    equaln #(12) e3072(.a(buffered_input), .b(12'b110000000000), .eq(weq3072));
    equaln #(12) e3073(.a(buffered_input), .b(12'b110000000001), .eq(weq3073));
    equaln #(12) e3074(.a(buffered_input), .b(12'b110000000010), .eq(weq3074));
    equaln #(12) e3075(.a(buffered_input), .b(12'b110000000011), .eq(weq3075));
    equaln #(12) e3076(.a(buffered_input), .b(12'b110000000100), .eq(weq3076));
    equaln #(12) e3077(.a(buffered_input), .b(12'b110000000101), .eq(weq3077));
    equaln #(12) e3078(.a(buffered_input), .b(12'b110000000110), .eq(weq3078));
    equaln #(12) e3079(.a(buffered_input), .b(12'b110000000111), .eq(weq3079));
    equaln #(12) e3080(.a(buffered_input), .b(12'b110000001000), .eq(weq3080));
    equaln #(12) e3081(.a(buffered_input), .b(12'b110000001001), .eq(weq3081));
    equaln #(12) e3082(.a(buffered_input), .b(12'b110000001010), .eq(weq3082));
    equaln #(12) e3083(.a(buffered_input), .b(12'b110000001011), .eq(weq3083));
    equaln #(12) e3084(.a(buffered_input), .b(12'b110000001100), .eq(weq3084));
    equaln #(12) e3085(.a(buffered_input), .b(12'b110000001101), .eq(weq3085));
    equaln #(12) e3086(.a(buffered_input), .b(12'b110000001110), .eq(weq3086));
    equaln #(12) e3087(.a(buffered_input), .b(12'b110000001111), .eq(weq3087));
    equaln #(12) e3088(.a(buffered_input), .b(12'b110000010000), .eq(weq3088));
    equaln #(12) e3089(.a(buffered_input), .b(12'b110000010001), .eq(weq3089));
    equaln #(12) e3090(.a(buffered_input), .b(12'b110000010010), .eq(weq3090));
    equaln #(12) e3091(.a(buffered_input), .b(12'b110000010011), .eq(weq3091));
    equaln #(12) e3092(.a(buffered_input), .b(12'b110000010100), .eq(weq3092));
    equaln #(12) e3093(.a(buffered_input), .b(12'b110000010101), .eq(weq3093));
    equaln #(12) e3094(.a(buffered_input), .b(12'b110000010110), .eq(weq3094));
    equaln #(12) e3095(.a(buffered_input), .b(12'b110000010111), .eq(weq3095));
    equaln #(12) e3096(.a(buffered_input), .b(12'b110000011000), .eq(weq3096));
    equaln #(12) e3097(.a(buffered_input), .b(12'b110000011001), .eq(weq3097));
    equaln #(12) e3098(.a(buffered_input), .b(12'b110000011010), .eq(weq3098));
    equaln #(12) e3099(.a(buffered_input), .b(12'b110000011011), .eq(weq3099));
    equaln #(12) e3100(.a(buffered_input), .b(12'b110000011100), .eq(weq3100));
    equaln #(12) e3101(.a(buffered_input), .b(12'b110000011101), .eq(weq3101));
    equaln #(12) e3102(.a(buffered_input), .b(12'b110000011110), .eq(weq3102));
    equaln #(12) e3103(.a(buffered_input), .b(12'b110000011111), .eq(weq3103));
    equaln #(12) e3104(.a(buffered_input), .b(12'b110000100000), .eq(weq3104));
    equaln #(12) e3105(.a(buffered_input), .b(12'b110000100001), .eq(weq3105));
    equaln #(12) e3106(.a(buffered_input), .b(12'b110000100010), .eq(weq3106));
    equaln #(12) e3107(.a(buffered_input), .b(12'b110000100011), .eq(weq3107));
    equaln #(12) e3108(.a(buffered_input), .b(12'b110000100100), .eq(weq3108));
    equaln #(12) e3109(.a(buffered_input), .b(12'b110000100101), .eq(weq3109));
    equaln #(12) e3110(.a(buffered_input), .b(12'b110000100110), .eq(weq3110));
    equaln #(12) e3111(.a(buffered_input), .b(12'b110000100111), .eq(weq3111));
    equaln #(12) e3112(.a(buffered_input), .b(12'b110000101000), .eq(weq3112));
    equaln #(12) e3113(.a(buffered_input), .b(12'b110000101001), .eq(weq3113));
    equaln #(12) e3114(.a(buffered_input), .b(12'b110000101010), .eq(weq3114));
    equaln #(12) e3115(.a(buffered_input), .b(12'b110000101011), .eq(weq3115));
    equaln #(12) e3116(.a(buffered_input), .b(12'b110000101100), .eq(weq3116));
    equaln #(12) e3117(.a(buffered_input), .b(12'b110000101101), .eq(weq3117));
    equaln #(12) e3118(.a(buffered_input), .b(12'b110000101110), .eq(weq3118));
    equaln #(12) e3119(.a(buffered_input), .b(12'b110000101111), .eq(weq3119));
    equaln #(12) e3120(.a(buffered_input), .b(12'b110000110000), .eq(weq3120));
    equaln #(12) e3121(.a(buffered_input), .b(12'b110000110001), .eq(weq3121));
    equaln #(12) e3122(.a(buffered_input), .b(12'b110000110010), .eq(weq3122));
    equaln #(12) e3123(.a(buffered_input), .b(12'b110000110011), .eq(weq3123));
    equaln #(12) e3124(.a(buffered_input), .b(12'b110000110100), .eq(weq3124));
    equaln #(12) e3125(.a(buffered_input), .b(12'b110000110101), .eq(weq3125));
    equaln #(12) e3126(.a(buffered_input), .b(12'b110000110110), .eq(weq3126));
    equaln #(12) e3127(.a(buffered_input), .b(12'b110000110111), .eq(weq3127));
    equaln #(12) e3128(.a(buffered_input), .b(12'b110000111000), .eq(weq3128));
    equaln #(12) e3129(.a(buffered_input), .b(12'b110000111001), .eq(weq3129));
    equaln #(12) e3130(.a(buffered_input), .b(12'b110000111010), .eq(weq3130));
    equaln #(12) e3131(.a(buffered_input), .b(12'b110000111011), .eq(weq3131));
    equaln #(12) e3132(.a(buffered_input), .b(12'b110000111100), .eq(weq3132));
    equaln #(12) e3133(.a(buffered_input), .b(12'b110000111101), .eq(weq3133));
    equaln #(12) e3134(.a(buffered_input), .b(12'b110000111110), .eq(weq3134));
    equaln #(12) e3135(.a(buffered_input), .b(12'b110000111111), .eq(weq3135));
    equaln #(12) e3136(.a(buffered_input), .b(12'b110001000000), .eq(weq3136));
    equaln #(12) e3137(.a(buffered_input), .b(12'b110001000001), .eq(weq3137));
    equaln #(12) e3138(.a(buffered_input), .b(12'b110001000010), .eq(weq3138));
    equaln #(12) e3139(.a(buffered_input), .b(12'b110001000011), .eq(weq3139));
    equaln #(12) e3140(.a(buffered_input), .b(12'b110001000100), .eq(weq3140));
    equaln #(12) e3141(.a(buffered_input), .b(12'b110001000101), .eq(weq3141));
    equaln #(12) e3142(.a(buffered_input), .b(12'b110001000110), .eq(weq3142));
    equaln #(12) e3143(.a(buffered_input), .b(12'b110001000111), .eq(weq3143));
    equaln #(12) e3144(.a(buffered_input), .b(12'b110001001000), .eq(weq3144));
    equaln #(12) e3145(.a(buffered_input), .b(12'b110001001001), .eq(weq3145));
    equaln #(12) e3146(.a(buffered_input), .b(12'b110001001010), .eq(weq3146));
    equaln #(12) e3147(.a(buffered_input), .b(12'b110001001011), .eq(weq3147));
    equaln #(12) e3148(.a(buffered_input), .b(12'b110001001100), .eq(weq3148));
    equaln #(12) e3149(.a(buffered_input), .b(12'b110001001101), .eq(weq3149));
    equaln #(12) e3150(.a(buffered_input), .b(12'b110001001110), .eq(weq3150));
    equaln #(12) e3151(.a(buffered_input), .b(12'b110001001111), .eq(weq3151));
    equaln #(12) e3152(.a(buffered_input), .b(12'b110001010000), .eq(weq3152));
    equaln #(12) e3153(.a(buffered_input), .b(12'b110001010001), .eq(weq3153));
    equaln #(12) e3154(.a(buffered_input), .b(12'b110001010010), .eq(weq3154));
    equaln #(12) e3155(.a(buffered_input), .b(12'b110001010011), .eq(weq3155));
    equaln #(12) e3156(.a(buffered_input), .b(12'b110001010100), .eq(weq3156));
    equaln #(12) e3157(.a(buffered_input), .b(12'b110001010101), .eq(weq3157));
    equaln #(12) e3158(.a(buffered_input), .b(12'b110001010110), .eq(weq3158));
    equaln #(12) e3159(.a(buffered_input), .b(12'b110001010111), .eq(weq3159));
    equaln #(12) e3160(.a(buffered_input), .b(12'b110001011000), .eq(weq3160));
    equaln #(12) e3161(.a(buffered_input), .b(12'b110001011001), .eq(weq3161));
    equaln #(12) e3162(.a(buffered_input), .b(12'b110001011010), .eq(weq3162));
    equaln #(12) e3163(.a(buffered_input), .b(12'b110001011011), .eq(weq3163));
    equaln #(12) e3164(.a(buffered_input), .b(12'b110001011100), .eq(weq3164));
    equaln #(12) e3165(.a(buffered_input), .b(12'b110001011101), .eq(weq3165));
    equaln #(12) e3166(.a(buffered_input), .b(12'b110001011110), .eq(weq3166));
    equaln #(12) e3167(.a(buffered_input), .b(12'b110001011111), .eq(weq3167));
    equaln #(12) e3168(.a(buffered_input), .b(12'b110001100000), .eq(weq3168));
    equaln #(12) e3169(.a(buffered_input), .b(12'b110001100001), .eq(weq3169));
    equaln #(12) e3170(.a(buffered_input), .b(12'b110001100010), .eq(weq3170));
    equaln #(12) e3171(.a(buffered_input), .b(12'b110001100011), .eq(weq3171));
    equaln #(12) e3172(.a(buffered_input), .b(12'b110001100100), .eq(weq3172));
    equaln #(12) e3173(.a(buffered_input), .b(12'b110001100101), .eq(weq3173));
    equaln #(12) e3174(.a(buffered_input), .b(12'b110001100110), .eq(weq3174));
    equaln #(12) e3175(.a(buffered_input), .b(12'b110001100111), .eq(weq3175));
    equaln #(12) e3176(.a(buffered_input), .b(12'b110001101000), .eq(weq3176));
    equaln #(12) e3177(.a(buffered_input), .b(12'b110001101001), .eq(weq3177));
    equaln #(12) e3178(.a(buffered_input), .b(12'b110001101010), .eq(weq3178));
    equaln #(12) e3179(.a(buffered_input), .b(12'b110001101011), .eq(weq3179));
    equaln #(12) e3180(.a(buffered_input), .b(12'b110001101100), .eq(weq3180));
    equaln #(12) e3181(.a(buffered_input), .b(12'b110001101101), .eq(weq3181));
    equaln #(12) e3182(.a(buffered_input), .b(12'b110001101110), .eq(weq3182));
    equaln #(12) e3183(.a(buffered_input), .b(12'b110001101111), .eq(weq3183));
    equaln #(12) e3184(.a(buffered_input), .b(12'b110001110000), .eq(weq3184));
    equaln #(12) e3185(.a(buffered_input), .b(12'b110001110001), .eq(weq3185));
    equaln #(12) e3186(.a(buffered_input), .b(12'b110001110010), .eq(weq3186));
    equaln #(12) e3187(.a(buffered_input), .b(12'b110001110011), .eq(weq3187));
    equaln #(12) e3188(.a(buffered_input), .b(12'b110001110100), .eq(weq3188));
    equaln #(12) e3189(.a(buffered_input), .b(12'b110001110101), .eq(weq3189));
    equaln #(12) e3190(.a(buffered_input), .b(12'b110001110110), .eq(weq3190));
    equaln #(12) e3191(.a(buffered_input), .b(12'b110001110111), .eq(weq3191));
    equaln #(12) e3192(.a(buffered_input), .b(12'b110001111000), .eq(weq3192));
    equaln #(12) e3193(.a(buffered_input), .b(12'b110001111001), .eq(weq3193));
    equaln #(12) e3194(.a(buffered_input), .b(12'b110001111010), .eq(weq3194));
    equaln #(12) e3195(.a(buffered_input), .b(12'b110001111011), .eq(weq3195));
    equaln #(12) e3196(.a(buffered_input), .b(12'b110001111100), .eq(weq3196));
    equaln #(12) e3197(.a(buffered_input), .b(12'b110001111101), .eq(weq3197));
    equaln #(12) e3198(.a(buffered_input), .b(12'b110001111110), .eq(weq3198));
    equaln #(12) e3199(.a(buffered_input), .b(12'b110001111111), .eq(weq3199));
    equaln #(12) e3200(.a(buffered_input), .b(12'b110010000000), .eq(weq3200));
    equaln #(12) e3201(.a(buffered_input), .b(12'b110010000001), .eq(weq3201));
    equaln #(12) e3202(.a(buffered_input), .b(12'b110010000010), .eq(weq3202));
    equaln #(12) e3203(.a(buffered_input), .b(12'b110010000011), .eq(weq3203));
    equaln #(12) e3204(.a(buffered_input), .b(12'b110010000100), .eq(weq3204));
    equaln #(12) e3205(.a(buffered_input), .b(12'b110010000101), .eq(weq3205));
    equaln #(12) e3206(.a(buffered_input), .b(12'b110010000110), .eq(weq3206));
    equaln #(12) e3207(.a(buffered_input), .b(12'b110010000111), .eq(weq3207));
    equaln #(12) e3208(.a(buffered_input), .b(12'b110010001000), .eq(weq3208));
    equaln #(12) e3209(.a(buffered_input), .b(12'b110010001001), .eq(weq3209));
    equaln #(12) e3210(.a(buffered_input), .b(12'b110010001010), .eq(weq3210));
    equaln #(12) e3211(.a(buffered_input), .b(12'b110010001011), .eq(weq3211));
    equaln #(12) e3212(.a(buffered_input), .b(12'b110010001100), .eq(weq3212));
    equaln #(12) e3213(.a(buffered_input), .b(12'b110010001101), .eq(weq3213));
    equaln #(12) e3214(.a(buffered_input), .b(12'b110010001110), .eq(weq3214));
    equaln #(12) e3215(.a(buffered_input), .b(12'b110010001111), .eq(weq3215));
    equaln #(12) e3216(.a(buffered_input), .b(12'b110010010000), .eq(weq3216));
    equaln #(12) e3217(.a(buffered_input), .b(12'b110010010001), .eq(weq3217));
    equaln #(12) e3218(.a(buffered_input), .b(12'b110010010010), .eq(weq3218));
    equaln #(12) e3219(.a(buffered_input), .b(12'b110010010011), .eq(weq3219));
    equaln #(12) e3220(.a(buffered_input), .b(12'b110010010100), .eq(weq3220));
    equaln #(12) e3221(.a(buffered_input), .b(12'b110010010101), .eq(weq3221));
    equaln #(12) e3222(.a(buffered_input), .b(12'b110010010110), .eq(weq3222));
    equaln #(12) e3223(.a(buffered_input), .b(12'b110010010111), .eq(weq3223));
    equaln #(12) e3224(.a(buffered_input), .b(12'b110010011000), .eq(weq3224));
    equaln #(12) e3225(.a(buffered_input), .b(12'b110010011001), .eq(weq3225));
    equaln #(12) e3226(.a(buffered_input), .b(12'b110010011010), .eq(weq3226));
    equaln #(12) e3227(.a(buffered_input), .b(12'b110010011011), .eq(weq3227));
    equaln #(12) e3228(.a(buffered_input), .b(12'b110010011100), .eq(weq3228));
    equaln #(12) e3229(.a(buffered_input), .b(12'b110010011101), .eq(weq3229));
    equaln #(12) e3230(.a(buffered_input), .b(12'b110010011110), .eq(weq3230));
    equaln #(12) e3231(.a(buffered_input), .b(12'b110010011111), .eq(weq3231));
    equaln #(12) e3232(.a(buffered_input), .b(12'b110010100000), .eq(weq3232));
    equaln #(12) e3233(.a(buffered_input), .b(12'b110010100001), .eq(weq3233));
    equaln #(12) e3234(.a(buffered_input), .b(12'b110010100010), .eq(weq3234));
    equaln #(12) e3235(.a(buffered_input), .b(12'b110010100011), .eq(weq3235));
    equaln #(12) e3236(.a(buffered_input), .b(12'b110010100100), .eq(weq3236));
    equaln #(12) e3237(.a(buffered_input), .b(12'b110010100101), .eq(weq3237));
    equaln #(12) e3238(.a(buffered_input), .b(12'b110010100110), .eq(weq3238));
    equaln #(12) e3239(.a(buffered_input), .b(12'b110010100111), .eq(weq3239));
    equaln #(12) e3240(.a(buffered_input), .b(12'b110010101000), .eq(weq3240));
    equaln #(12) e3241(.a(buffered_input), .b(12'b110010101001), .eq(weq3241));
    equaln #(12) e3242(.a(buffered_input), .b(12'b110010101010), .eq(weq3242));
    equaln #(12) e3243(.a(buffered_input), .b(12'b110010101011), .eq(weq3243));
    equaln #(12) e3244(.a(buffered_input), .b(12'b110010101100), .eq(weq3244));
    equaln #(12) e3245(.a(buffered_input), .b(12'b110010101101), .eq(weq3245));
    equaln #(12) e3246(.a(buffered_input), .b(12'b110010101110), .eq(weq3246));
    equaln #(12) e3247(.a(buffered_input), .b(12'b110010101111), .eq(weq3247));
    equaln #(12) e3248(.a(buffered_input), .b(12'b110010110000), .eq(weq3248));
    equaln #(12) e3249(.a(buffered_input), .b(12'b110010110001), .eq(weq3249));
    equaln #(12) e3250(.a(buffered_input), .b(12'b110010110010), .eq(weq3250));
    equaln #(12) e3251(.a(buffered_input), .b(12'b110010110011), .eq(weq3251));
    equaln #(12) e3252(.a(buffered_input), .b(12'b110010110100), .eq(weq3252));
    equaln #(12) e3253(.a(buffered_input), .b(12'b110010110101), .eq(weq3253));
    equaln #(12) e3254(.a(buffered_input), .b(12'b110010110110), .eq(weq3254));
    equaln #(12) e3255(.a(buffered_input), .b(12'b110010110111), .eq(weq3255));
    equaln #(12) e3256(.a(buffered_input), .b(12'b110010111000), .eq(weq3256));
    equaln #(12) e3257(.a(buffered_input), .b(12'b110010111001), .eq(weq3257));
    equaln #(12) e3258(.a(buffered_input), .b(12'b110010111010), .eq(weq3258));
    equaln #(12) e3259(.a(buffered_input), .b(12'b110010111011), .eq(weq3259));
    equaln #(12) e3260(.a(buffered_input), .b(12'b110010111100), .eq(weq3260));
    equaln #(12) e3261(.a(buffered_input), .b(12'b110010111101), .eq(weq3261));
    equaln #(12) e3262(.a(buffered_input), .b(12'b110010111110), .eq(weq3262));
    equaln #(12) e3263(.a(buffered_input), .b(12'b110010111111), .eq(weq3263));
    equaln #(12) e3264(.a(buffered_input), .b(12'b110011000000), .eq(weq3264));
    equaln #(12) e3265(.a(buffered_input), .b(12'b110011000001), .eq(weq3265));
    equaln #(12) e3266(.a(buffered_input), .b(12'b110011000010), .eq(weq3266));
    equaln #(12) e3267(.a(buffered_input), .b(12'b110011000011), .eq(weq3267));
    equaln #(12) e3268(.a(buffered_input), .b(12'b110011000100), .eq(weq3268));
    equaln #(12) e3269(.a(buffered_input), .b(12'b110011000101), .eq(weq3269));
    equaln #(12) e3270(.a(buffered_input), .b(12'b110011000110), .eq(weq3270));
    equaln #(12) e3271(.a(buffered_input), .b(12'b110011000111), .eq(weq3271));
    equaln #(12) e3272(.a(buffered_input), .b(12'b110011001000), .eq(weq3272));
    equaln #(12) e3273(.a(buffered_input), .b(12'b110011001001), .eq(weq3273));
    equaln #(12) e3274(.a(buffered_input), .b(12'b110011001010), .eq(weq3274));
    equaln #(12) e3275(.a(buffered_input), .b(12'b110011001011), .eq(weq3275));
    equaln #(12) e3276(.a(buffered_input), .b(12'b110011001100), .eq(weq3276));
    equaln #(12) e3277(.a(buffered_input), .b(12'b110011001101), .eq(weq3277));
    equaln #(12) e3278(.a(buffered_input), .b(12'b110011001110), .eq(weq3278));
    equaln #(12) e3279(.a(buffered_input), .b(12'b110011001111), .eq(weq3279));
    equaln #(12) e3280(.a(buffered_input), .b(12'b110011010000), .eq(weq3280));
    equaln #(12) e3281(.a(buffered_input), .b(12'b110011010001), .eq(weq3281));
    equaln #(12) e3282(.a(buffered_input), .b(12'b110011010010), .eq(weq3282));
    equaln #(12) e3283(.a(buffered_input), .b(12'b110011010011), .eq(weq3283));
    equaln #(12) e3284(.a(buffered_input), .b(12'b110011010100), .eq(weq3284));
    equaln #(12) e3285(.a(buffered_input), .b(12'b110011010101), .eq(weq3285));
    equaln #(12) e3286(.a(buffered_input), .b(12'b110011010110), .eq(weq3286));
    equaln #(12) e3287(.a(buffered_input), .b(12'b110011010111), .eq(weq3287));
    equaln #(12) e3288(.a(buffered_input), .b(12'b110011011000), .eq(weq3288));
    equaln #(12) e3289(.a(buffered_input), .b(12'b110011011001), .eq(weq3289));
    equaln #(12) e3290(.a(buffered_input), .b(12'b110011011010), .eq(weq3290));
    equaln #(12) e3291(.a(buffered_input), .b(12'b110011011011), .eq(weq3291));
    equaln #(12) e3292(.a(buffered_input), .b(12'b110011011100), .eq(weq3292));
    equaln #(12) e3293(.a(buffered_input), .b(12'b110011011101), .eq(weq3293));
    equaln #(12) e3294(.a(buffered_input), .b(12'b110011011110), .eq(weq3294));
    equaln #(12) e3295(.a(buffered_input), .b(12'b110011011111), .eq(weq3295));
    equaln #(12) e3296(.a(buffered_input), .b(12'b110011100000), .eq(weq3296));
    equaln #(12) e3297(.a(buffered_input), .b(12'b110011100001), .eq(weq3297));
    equaln #(12) e3298(.a(buffered_input), .b(12'b110011100010), .eq(weq3298));
    equaln #(12) e3299(.a(buffered_input), .b(12'b110011100011), .eq(weq3299));
    equaln #(12) e3300(.a(buffered_input), .b(12'b110011100100), .eq(weq3300));
    equaln #(12) e3301(.a(buffered_input), .b(12'b110011100101), .eq(weq3301));
    equaln #(12) e3302(.a(buffered_input), .b(12'b110011100110), .eq(weq3302));
    equaln #(12) e3303(.a(buffered_input), .b(12'b110011100111), .eq(weq3303));
    equaln #(12) e3304(.a(buffered_input), .b(12'b110011101000), .eq(weq3304));
    equaln #(12) e3305(.a(buffered_input), .b(12'b110011101001), .eq(weq3305));
    equaln #(12) e3306(.a(buffered_input), .b(12'b110011101010), .eq(weq3306));
    equaln #(12) e3307(.a(buffered_input), .b(12'b110011101011), .eq(weq3307));
    equaln #(12) e3308(.a(buffered_input), .b(12'b110011101100), .eq(weq3308));
    equaln #(12) e3309(.a(buffered_input), .b(12'b110011101101), .eq(weq3309));
    equaln #(12) e3310(.a(buffered_input), .b(12'b110011101110), .eq(weq3310));
    equaln #(12) e3311(.a(buffered_input), .b(12'b110011101111), .eq(weq3311));
    equaln #(12) e3312(.a(buffered_input), .b(12'b110011110000), .eq(weq3312));
    equaln #(12) e3313(.a(buffered_input), .b(12'b110011110001), .eq(weq3313));
    equaln #(12) e3314(.a(buffered_input), .b(12'b110011110010), .eq(weq3314));
    equaln #(12) e3315(.a(buffered_input), .b(12'b110011110011), .eq(weq3315));
    equaln #(12) e3316(.a(buffered_input), .b(12'b110011110100), .eq(weq3316));
    equaln #(12) e3317(.a(buffered_input), .b(12'b110011110101), .eq(weq3317));
    equaln #(12) e3318(.a(buffered_input), .b(12'b110011110110), .eq(weq3318));
    equaln #(12) e3319(.a(buffered_input), .b(12'b110011110111), .eq(weq3319));
    equaln #(12) e3320(.a(buffered_input), .b(12'b110011111000), .eq(weq3320));
    equaln #(12) e3321(.a(buffered_input), .b(12'b110011111001), .eq(weq3321));
    equaln #(12) e3322(.a(buffered_input), .b(12'b110011111010), .eq(weq3322));
    equaln #(12) e3323(.a(buffered_input), .b(12'b110011111011), .eq(weq3323));
    equaln #(12) e3324(.a(buffered_input), .b(12'b110011111100), .eq(weq3324));
    equaln #(12) e3325(.a(buffered_input), .b(12'b110011111101), .eq(weq3325));
    equaln #(12) e3326(.a(buffered_input), .b(12'b110011111110), .eq(weq3326));
    equaln #(12) e3327(.a(buffered_input), .b(12'b110011111111), .eq(weq3327));
    equaln #(12) e3328(.a(buffered_input), .b(12'b110100000000), .eq(weq3328));
    equaln #(12) e3329(.a(buffered_input), .b(12'b110100000001), .eq(weq3329));
    equaln #(12) e3330(.a(buffered_input), .b(12'b110100000010), .eq(weq3330));
    equaln #(12) e3331(.a(buffered_input), .b(12'b110100000011), .eq(weq3331));
    equaln #(12) e3332(.a(buffered_input), .b(12'b110100000100), .eq(weq3332));
    equaln #(12) e3333(.a(buffered_input), .b(12'b110100000101), .eq(weq3333));
    equaln #(12) e3334(.a(buffered_input), .b(12'b110100000110), .eq(weq3334));
    equaln #(12) e3335(.a(buffered_input), .b(12'b110100000111), .eq(weq3335));
    equaln #(12) e3336(.a(buffered_input), .b(12'b110100001000), .eq(weq3336));
    equaln #(12) e3337(.a(buffered_input), .b(12'b110100001001), .eq(weq3337));
    equaln #(12) e3338(.a(buffered_input), .b(12'b110100001010), .eq(weq3338));
    equaln #(12) e3339(.a(buffered_input), .b(12'b110100001011), .eq(weq3339));
    equaln #(12) e3340(.a(buffered_input), .b(12'b110100001100), .eq(weq3340));
    equaln #(12) e3341(.a(buffered_input), .b(12'b110100001101), .eq(weq3341));
    equaln #(12) e3342(.a(buffered_input), .b(12'b110100001110), .eq(weq3342));
    equaln #(12) e3343(.a(buffered_input), .b(12'b110100001111), .eq(weq3343));
    equaln #(12) e3344(.a(buffered_input), .b(12'b110100010000), .eq(weq3344));
    equaln #(12) e3345(.a(buffered_input), .b(12'b110100010001), .eq(weq3345));
    equaln #(12) e3346(.a(buffered_input), .b(12'b110100010010), .eq(weq3346));
    equaln #(12) e3347(.a(buffered_input), .b(12'b110100010011), .eq(weq3347));
    equaln #(12) e3348(.a(buffered_input), .b(12'b110100010100), .eq(weq3348));
    equaln #(12) e3349(.a(buffered_input), .b(12'b110100010101), .eq(weq3349));
    equaln #(12) e3350(.a(buffered_input), .b(12'b110100010110), .eq(weq3350));
    equaln #(12) e3351(.a(buffered_input), .b(12'b110100010111), .eq(weq3351));
    equaln #(12) e3352(.a(buffered_input), .b(12'b110100011000), .eq(weq3352));
    equaln #(12) e3353(.a(buffered_input), .b(12'b110100011001), .eq(weq3353));
    equaln #(12) e3354(.a(buffered_input), .b(12'b110100011010), .eq(weq3354));
    equaln #(12) e3355(.a(buffered_input), .b(12'b110100011011), .eq(weq3355));
    equaln #(12) e3356(.a(buffered_input), .b(12'b110100011100), .eq(weq3356));
    equaln #(12) e3357(.a(buffered_input), .b(12'b110100011101), .eq(weq3357));
    equaln #(12) e3358(.a(buffered_input), .b(12'b110100011110), .eq(weq3358));
    equaln #(12) e3359(.a(buffered_input), .b(12'b110100011111), .eq(weq3359));
    equaln #(12) e3360(.a(buffered_input), .b(12'b110100100000), .eq(weq3360));
    equaln #(12) e3361(.a(buffered_input), .b(12'b110100100001), .eq(weq3361));
    equaln #(12) e3362(.a(buffered_input), .b(12'b110100100010), .eq(weq3362));
    equaln #(12) e3363(.a(buffered_input), .b(12'b110100100011), .eq(weq3363));
    equaln #(12) e3364(.a(buffered_input), .b(12'b110100100100), .eq(weq3364));
    equaln #(12) e3365(.a(buffered_input), .b(12'b110100100101), .eq(weq3365));
    equaln #(12) e3366(.a(buffered_input), .b(12'b110100100110), .eq(weq3366));
    equaln #(12) e3367(.a(buffered_input), .b(12'b110100100111), .eq(weq3367));
    equaln #(12) e3368(.a(buffered_input), .b(12'b110100101000), .eq(weq3368));
    equaln #(12) e3369(.a(buffered_input), .b(12'b110100101001), .eq(weq3369));
    equaln #(12) e3370(.a(buffered_input), .b(12'b110100101010), .eq(weq3370));
    equaln #(12) e3371(.a(buffered_input), .b(12'b110100101011), .eq(weq3371));
    equaln #(12) e3372(.a(buffered_input), .b(12'b110100101100), .eq(weq3372));
    equaln #(12) e3373(.a(buffered_input), .b(12'b110100101101), .eq(weq3373));
    equaln #(12) e3374(.a(buffered_input), .b(12'b110100101110), .eq(weq3374));
    equaln #(12) e3375(.a(buffered_input), .b(12'b110100101111), .eq(weq3375));
    equaln #(12) e3376(.a(buffered_input), .b(12'b110100110000), .eq(weq3376));
    equaln #(12) e3377(.a(buffered_input), .b(12'b110100110001), .eq(weq3377));
    equaln #(12) e3378(.a(buffered_input), .b(12'b110100110010), .eq(weq3378));
    equaln #(12) e3379(.a(buffered_input), .b(12'b110100110011), .eq(weq3379));
    equaln #(12) e3380(.a(buffered_input), .b(12'b110100110100), .eq(weq3380));
    equaln #(12) e3381(.a(buffered_input), .b(12'b110100110101), .eq(weq3381));
    equaln #(12) e3382(.a(buffered_input), .b(12'b110100110110), .eq(weq3382));
    equaln #(12) e3383(.a(buffered_input), .b(12'b110100110111), .eq(weq3383));
    equaln #(12) e3384(.a(buffered_input), .b(12'b110100111000), .eq(weq3384));
    equaln #(12) e3385(.a(buffered_input), .b(12'b110100111001), .eq(weq3385));
    equaln #(12) e3386(.a(buffered_input), .b(12'b110100111010), .eq(weq3386));
    equaln #(12) e3387(.a(buffered_input), .b(12'b110100111011), .eq(weq3387));
    equaln #(12) e3388(.a(buffered_input), .b(12'b110100111100), .eq(weq3388));
    equaln #(12) e3389(.a(buffered_input), .b(12'b110100111101), .eq(weq3389));
    equaln #(12) e3390(.a(buffered_input), .b(12'b110100111110), .eq(weq3390));
    equaln #(12) e3391(.a(buffered_input), .b(12'b110100111111), .eq(weq3391));
    equaln #(12) e3392(.a(buffered_input), .b(12'b110101000000), .eq(weq3392));
    equaln #(12) e3393(.a(buffered_input), .b(12'b110101000001), .eq(weq3393));
    equaln #(12) e3394(.a(buffered_input), .b(12'b110101000010), .eq(weq3394));
    equaln #(12) e3395(.a(buffered_input), .b(12'b110101000011), .eq(weq3395));
    equaln #(12) e3396(.a(buffered_input), .b(12'b110101000100), .eq(weq3396));
    equaln #(12) e3397(.a(buffered_input), .b(12'b110101000101), .eq(weq3397));
    equaln #(12) e3398(.a(buffered_input), .b(12'b110101000110), .eq(weq3398));
    equaln #(12) e3399(.a(buffered_input), .b(12'b110101000111), .eq(weq3399));
    equaln #(12) e3400(.a(buffered_input), .b(12'b110101001000), .eq(weq3400));
    equaln #(12) e3401(.a(buffered_input), .b(12'b110101001001), .eq(weq3401));
    equaln #(12) e3402(.a(buffered_input), .b(12'b110101001010), .eq(weq3402));
    equaln #(12) e3403(.a(buffered_input), .b(12'b110101001011), .eq(weq3403));
    equaln #(12) e3404(.a(buffered_input), .b(12'b110101001100), .eq(weq3404));
    equaln #(12) e3405(.a(buffered_input), .b(12'b110101001101), .eq(weq3405));
    equaln #(12) e3406(.a(buffered_input), .b(12'b110101001110), .eq(weq3406));
    equaln #(12) e3407(.a(buffered_input), .b(12'b110101001111), .eq(weq3407));
    equaln #(12) e3408(.a(buffered_input), .b(12'b110101010000), .eq(weq3408));
    equaln #(12) e3409(.a(buffered_input), .b(12'b110101010001), .eq(weq3409));
    equaln #(12) e3410(.a(buffered_input), .b(12'b110101010010), .eq(weq3410));
    equaln #(12) e3411(.a(buffered_input), .b(12'b110101010011), .eq(weq3411));
    equaln #(12) e3412(.a(buffered_input), .b(12'b110101010100), .eq(weq3412));
    equaln #(12) e3413(.a(buffered_input), .b(12'b110101010101), .eq(weq3413));
    equaln #(12) e3414(.a(buffered_input), .b(12'b110101010110), .eq(weq3414));
    equaln #(12) e3415(.a(buffered_input), .b(12'b110101010111), .eq(weq3415));
    equaln #(12) e3416(.a(buffered_input), .b(12'b110101011000), .eq(weq3416));
    equaln #(12) e3417(.a(buffered_input), .b(12'b110101011001), .eq(weq3417));
    equaln #(12) e3418(.a(buffered_input), .b(12'b110101011010), .eq(weq3418));
    equaln #(12) e3419(.a(buffered_input), .b(12'b110101011011), .eq(weq3419));
    equaln #(12) e3420(.a(buffered_input), .b(12'b110101011100), .eq(weq3420));
    equaln #(12) e3421(.a(buffered_input), .b(12'b110101011101), .eq(weq3421));
    equaln #(12) e3422(.a(buffered_input), .b(12'b110101011110), .eq(weq3422));
    equaln #(12) e3423(.a(buffered_input), .b(12'b110101011111), .eq(weq3423));
    equaln #(12) e3424(.a(buffered_input), .b(12'b110101100000), .eq(weq3424));
    equaln #(12) e3425(.a(buffered_input), .b(12'b110101100001), .eq(weq3425));
    equaln #(12) e3426(.a(buffered_input), .b(12'b110101100010), .eq(weq3426));
    equaln #(12) e3427(.a(buffered_input), .b(12'b110101100011), .eq(weq3427));
    equaln #(12) e3428(.a(buffered_input), .b(12'b110101100100), .eq(weq3428));
    equaln #(12) e3429(.a(buffered_input), .b(12'b110101100101), .eq(weq3429));
    equaln #(12) e3430(.a(buffered_input), .b(12'b110101100110), .eq(weq3430));
    equaln #(12) e3431(.a(buffered_input), .b(12'b110101100111), .eq(weq3431));
    equaln #(12) e3432(.a(buffered_input), .b(12'b110101101000), .eq(weq3432));
    equaln #(12) e3433(.a(buffered_input), .b(12'b110101101001), .eq(weq3433));
    equaln #(12) e3434(.a(buffered_input), .b(12'b110101101010), .eq(weq3434));
    equaln #(12) e3435(.a(buffered_input), .b(12'b110101101011), .eq(weq3435));
    equaln #(12) e3436(.a(buffered_input), .b(12'b110101101100), .eq(weq3436));
    equaln #(12) e3437(.a(buffered_input), .b(12'b110101101101), .eq(weq3437));
    equaln #(12) e3438(.a(buffered_input), .b(12'b110101101110), .eq(weq3438));
    equaln #(12) e3439(.a(buffered_input), .b(12'b110101101111), .eq(weq3439));
    equaln #(12) e3440(.a(buffered_input), .b(12'b110101110000), .eq(weq3440));
    equaln #(12) e3441(.a(buffered_input), .b(12'b110101110001), .eq(weq3441));
    equaln #(12) e3442(.a(buffered_input), .b(12'b110101110010), .eq(weq3442));
    equaln #(12) e3443(.a(buffered_input), .b(12'b110101110011), .eq(weq3443));
    equaln #(12) e3444(.a(buffered_input), .b(12'b110101110100), .eq(weq3444));
    equaln #(12) e3445(.a(buffered_input), .b(12'b110101110101), .eq(weq3445));
    equaln #(12) e3446(.a(buffered_input), .b(12'b110101110110), .eq(weq3446));
    equaln #(12) e3447(.a(buffered_input), .b(12'b110101110111), .eq(weq3447));
    equaln #(12) e3448(.a(buffered_input), .b(12'b110101111000), .eq(weq3448));
    equaln #(12) e3449(.a(buffered_input), .b(12'b110101111001), .eq(weq3449));
    equaln #(12) e3450(.a(buffered_input), .b(12'b110101111010), .eq(weq3450));
    equaln #(12) e3451(.a(buffered_input), .b(12'b110101111011), .eq(weq3451));
    equaln #(12) e3452(.a(buffered_input), .b(12'b110101111100), .eq(weq3452));
    equaln #(12) e3453(.a(buffered_input), .b(12'b110101111101), .eq(weq3453));
    equaln #(12) e3454(.a(buffered_input), .b(12'b110101111110), .eq(weq3454));
    equaln #(12) e3455(.a(buffered_input), .b(12'b110101111111), .eq(weq3455));
    equaln #(12) e3456(.a(buffered_input), .b(12'b110110000000), .eq(weq3456));
    equaln #(12) e3457(.a(buffered_input), .b(12'b110110000001), .eq(weq3457));
    equaln #(12) e3458(.a(buffered_input), .b(12'b110110000010), .eq(weq3458));
    equaln #(12) e3459(.a(buffered_input), .b(12'b110110000011), .eq(weq3459));
    equaln #(12) e3460(.a(buffered_input), .b(12'b110110000100), .eq(weq3460));
    equaln #(12) e3461(.a(buffered_input), .b(12'b110110000101), .eq(weq3461));
    equaln #(12) e3462(.a(buffered_input), .b(12'b110110000110), .eq(weq3462));
    equaln #(12) e3463(.a(buffered_input), .b(12'b110110000111), .eq(weq3463));
    equaln #(12) e3464(.a(buffered_input), .b(12'b110110001000), .eq(weq3464));
    equaln #(12) e3465(.a(buffered_input), .b(12'b110110001001), .eq(weq3465));
    equaln #(12) e3466(.a(buffered_input), .b(12'b110110001010), .eq(weq3466));
    equaln #(12) e3467(.a(buffered_input), .b(12'b110110001011), .eq(weq3467));
    equaln #(12) e3468(.a(buffered_input), .b(12'b110110001100), .eq(weq3468));
    equaln #(12) e3469(.a(buffered_input), .b(12'b110110001101), .eq(weq3469));
    equaln #(12) e3470(.a(buffered_input), .b(12'b110110001110), .eq(weq3470));
    equaln #(12) e3471(.a(buffered_input), .b(12'b110110001111), .eq(weq3471));
    equaln #(12) e3472(.a(buffered_input), .b(12'b110110010000), .eq(weq3472));
    equaln #(12) e3473(.a(buffered_input), .b(12'b110110010001), .eq(weq3473));
    equaln #(12) e3474(.a(buffered_input), .b(12'b110110010010), .eq(weq3474));
    equaln #(12) e3475(.a(buffered_input), .b(12'b110110010011), .eq(weq3475));
    equaln #(12) e3476(.a(buffered_input), .b(12'b110110010100), .eq(weq3476));
    equaln #(12) e3477(.a(buffered_input), .b(12'b110110010101), .eq(weq3477));
    equaln #(12) e3478(.a(buffered_input), .b(12'b110110010110), .eq(weq3478));
    equaln #(12) e3479(.a(buffered_input), .b(12'b110110010111), .eq(weq3479));
    equaln #(12) e3480(.a(buffered_input), .b(12'b110110011000), .eq(weq3480));
    equaln #(12) e3481(.a(buffered_input), .b(12'b110110011001), .eq(weq3481));
    equaln #(12) e3482(.a(buffered_input), .b(12'b110110011010), .eq(weq3482));
    equaln #(12) e3483(.a(buffered_input), .b(12'b110110011011), .eq(weq3483));
    equaln #(12) e3484(.a(buffered_input), .b(12'b110110011100), .eq(weq3484));
    equaln #(12) e3485(.a(buffered_input), .b(12'b110110011101), .eq(weq3485));
    equaln #(12) e3486(.a(buffered_input), .b(12'b110110011110), .eq(weq3486));
    equaln #(12) e3487(.a(buffered_input), .b(12'b110110011111), .eq(weq3487));
    equaln #(12) e3488(.a(buffered_input), .b(12'b110110100000), .eq(weq3488));
    equaln #(12) e3489(.a(buffered_input), .b(12'b110110100001), .eq(weq3489));
    equaln #(12) e3490(.a(buffered_input), .b(12'b110110100010), .eq(weq3490));
    equaln #(12) e3491(.a(buffered_input), .b(12'b110110100011), .eq(weq3491));
    equaln #(12) e3492(.a(buffered_input), .b(12'b110110100100), .eq(weq3492));
    equaln #(12) e3493(.a(buffered_input), .b(12'b110110100101), .eq(weq3493));
    equaln #(12) e3494(.a(buffered_input), .b(12'b110110100110), .eq(weq3494));
    equaln #(12) e3495(.a(buffered_input), .b(12'b110110100111), .eq(weq3495));
    equaln #(12) e3496(.a(buffered_input), .b(12'b110110101000), .eq(weq3496));
    equaln #(12) e3497(.a(buffered_input), .b(12'b110110101001), .eq(weq3497));
    equaln #(12) e3498(.a(buffered_input), .b(12'b110110101010), .eq(weq3498));
    equaln #(12) e3499(.a(buffered_input), .b(12'b110110101011), .eq(weq3499));
    equaln #(12) e3500(.a(buffered_input), .b(12'b110110101100), .eq(weq3500));
    equaln #(12) e3501(.a(buffered_input), .b(12'b110110101101), .eq(weq3501));
    equaln #(12) e3502(.a(buffered_input), .b(12'b110110101110), .eq(weq3502));
    equaln #(12) e3503(.a(buffered_input), .b(12'b110110101111), .eq(weq3503));
    equaln #(12) e3504(.a(buffered_input), .b(12'b110110110000), .eq(weq3504));
    equaln #(12) e3505(.a(buffered_input), .b(12'b110110110001), .eq(weq3505));
    equaln #(12) e3506(.a(buffered_input), .b(12'b110110110010), .eq(weq3506));
    equaln #(12) e3507(.a(buffered_input), .b(12'b110110110011), .eq(weq3507));
    equaln #(12) e3508(.a(buffered_input), .b(12'b110110110100), .eq(weq3508));
    equaln #(12) e3509(.a(buffered_input), .b(12'b110110110101), .eq(weq3509));
    equaln #(12) e3510(.a(buffered_input), .b(12'b110110110110), .eq(weq3510));
    equaln #(12) e3511(.a(buffered_input), .b(12'b110110110111), .eq(weq3511));
    equaln #(12) e3512(.a(buffered_input), .b(12'b110110111000), .eq(weq3512));
    equaln #(12) e3513(.a(buffered_input), .b(12'b110110111001), .eq(weq3513));
    equaln #(12) e3514(.a(buffered_input), .b(12'b110110111010), .eq(weq3514));
    equaln #(12) e3515(.a(buffered_input), .b(12'b110110111011), .eq(weq3515));
    equaln #(12) e3516(.a(buffered_input), .b(12'b110110111100), .eq(weq3516));
    equaln #(12) e3517(.a(buffered_input), .b(12'b110110111101), .eq(weq3517));
    equaln #(12) e3518(.a(buffered_input), .b(12'b110110111110), .eq(weq3518));
    equaln #(12) e3519(.a(buffered_input), .b(12'b110110111111), .eq(weq3519));
    equaln #(12) e3520(.a(buffered_input), .b(12'b110111000000), .eq(weq3520));
    equaln #(12) e3521(.a(buffered_input), .b(12'b110111000001), .eq(weq3521));
    equaln #(12) e3522(.a(buffered_input), .b(12'b110111000010), .eq(weq3522));
    equaln #(12) e3523(.a(buffered_input), .b(12'b110111000011), .eq(weq3523));
    equaln #(12) e3524(.a(buffered_input), .b(12'b110111000100), .eq(weq3524));
    equaln #(12) e3525(.a(buffered_input), .b(12'b110111000101), .eq(weq3525));
    equaln #(12) e3526(.a(buffered_input), .b(12'b110111000110), .eq(weq3526));
    equaln #(12) e3527(.a(buffered_input), .b(12'b110111000111), .eq(weq3527));
    equaln #(12) e3528(.a(buffered_input), .b(12'b110111001000), .eq(weq3528));
    equaln #(12) e3529(.a(buffered_input), .b(12'b110111001001), .eq(weq3529));
    equaln #(12) e3530(.a(buffered_input), .b(12'b110111001010), .eq(weq3530));
    equaln #(12) e3531(.a(buffered_input), .b(12'b110111001011), .eq(weq3531));
    equaln #(12) e3532(.a(buffered_input), .b(12'b110111001100), .eq(weq3532));
    equaln #(12) e3533(.a(buffered_input), .b(12'b110111001101), .eq(weq3533));
    equaln #(12) e3534(.a(buffered_input), .b(12'b110111001110), .eq(weq3534));
    equaln #(12) e3535(.a(buffered_input), .b(12'b110111001111), .eq(weq3535));
    equaln #(12) e3536(.a(buffered_input), .b(12'b110111010000), .eq(weq3536));
    equaln #(12) e3537(.a(buffered_input), .b(12'b110111010001), .eq(weq3537));
    equaln #(12) e3538(.a(buffered_input), .b(12'b110111010010), .eq(weq3538));
    equaln #(12) e3539(.a(buffered_input), .b(12'b110111010011), .eq(weq3539));
    equaln #(12) e3540(.a(buffered_input), .b(12'b110111010100), .eq(weq3540));
    equaln #(12) e3541(.a(buffered_input), .b(12'b110111010101), .eq(weq3541));
    equaln #(12) e3542(.a(buffered_input), .b(12'b110111010110), .eq(weq3542));
    equaln #(12) e3543(.a(buffered_input), .b(12'b110111010111), .eq(weq3543));
    equaln #(12) e3544(.a(buffered_input), .b(12'b110111011000), .eq(weq3544));
    equaln #(12) e3545(.a(buffered_input), .b(12'b110111011001), .eq(weq3545));
    equaln #(12) e3546(.a(buffered_input), .b(12'b110111011010), .eq(weq3546));
    equaln #(12) e3547(.a(buffered_input), .b(12'b110111011011), .eq(weq3547));
    equaln #(12) e3548(.a(buffered_input), .b(12'b110111011100), .eq(weq3548));
    equaln #(12) e3549(.a(buffered_input), .b(12'b110111011101), .eq(weq3549));
    equaln #(12) e3550(.a(buffered_input), .b(12'b110111011110), .eq(weq3550));
    equaln #(12) e3551(.a(buffered_input), .b(12'b110111011111), .eq(weq3551));
    equaln #(12) e3552(.a(buffered_input), .b(12'b110111100000), .eq(weq3552));
    equaln #(12) e3553(.a(buffered_input), .b(12'b110111100001), .eq(weq3553));
    equaln #(12) e3554(.a(buffered_input), .b(12'b110111100010), .eq(weq3554));
    equaln #(12) e3555(.a(buffered_input), .b(12'b110111100011), .eq(weq3555));
    equaln #(12) e3556(.a(buffered_input), .b(12'b110111100100), .eq(weq3556));
    equaln #(12) e3557(.a(buffered_input), .b(12'b110111100101), .eq(weq3557));
    equaln #(12) e3558(.a(buffered_input), .b(12'b110111100110), .eq(weq3558));
    equaln #(12) e3559(.a(buffered_input), .b(12'b110111100111), .eq(weq3559));
    equaln #(12) e3560(.a(buffered_input), .b(12'b110111101000), .eq(weq3560));
    equaln #(12) e3561(.a(buffered_input), .b(12'b110111101001), .eq(weq3561));
    equaln #(12) e3562(.a(buffered_input), .b(12'b110111101010), .eq(weq3562));
    equaln #(12) e3563(.a(buffered_input), .b(12'b110111101011), .eq(weq3563));
    equaln #(12) e3564(.a(buffered_input), .b(12'b110111101100), .eq(weq3564));
    equaln #(12) e3565(.a(buffered_input), .b(12'b110111101101), .eq(weq3565));
    equaln #(12) e3566(.a(buffered_input), .b(12'b110111101110), .eq(weq3566));
    equaln #(12) e3567(.a(buffered_input), .b(12'b110111101111), .eq(weq3567));
    equaln #(12) e3568(.a(buffered_input), .b(12'b110111110000), .eq(weq3568));
    equaln #(12) e3569(.a(buffered_input), .b(12'b110111110001), .eq(weq3569));
    equaln #(12) e3570(.a(buffered_input), .b(12'b110111110010), .eq(weq3570));
    equaln #(12) e3571(.a(buffered_input), .b(12'b110111110011), .eq(weq3571));
    equaln #(12) e3572(.a(buffered_input), .b(12'b110111110100), .eq(weq3572));
    equaln #(12) e3573(.a(buffered_input), .b(12'b110111110101), .eq(weq3573));
    equaln #(12) e3574(.a(buffered_input), .b(12'b110111110110), .eq(weq3574));
    equaln #(12) e3575(.a(buffered_input), .b(12'b110111110111), .eq(weq3575));
    equaln #(12) e3576(.a(buffered_input), .b(12'b110111111000), .eq(weq3576));
    equaln #(12) e3577(.a(buffered_input), .b(12'b110111111001), .eq(weq3577));
    equaln #(12) e3578(.a(buffered_input), .b(12'b110111111010), .eq(weq3578));
    equaln #(12) e3579(.a(buffered_input), .b(12'b110111111011), .eq(weq3579));
    equaln #(12) e3580(.a(buffered_input), .b(12'b110111111100), .eq(weq3580));
    equaln #(12) e3581(.a(buffered_input), .b(12'b110111111101), .eq(weq3581));
    equaln #(12) e3582(.a(buffered_input), .b(12'b110111111110), .eq(weq3582));
    equaln #(12) e3583(.a(buffered_input), .b(12'b110111111111), .eq(weq3583));
    equaln #(12) e3584(.a(buffered_input), .b(12'b111000000000), .eq(weq3584));
    equaln #(12) e3585(.a(buffered_input), .b(12'b111000000001), .eq(weq3585));
    equaln #(12) e3586(.a(buffered_input), .b(12'b111000000010), .eq(weq3586));
    equaln #(12) e3587(.a(buffered_input), .b(12'b111000000011), .eq(weq3587));
    equaln #(12) e3588(.a(buffered_input), .b(12'b111000000100), .eq(weq3588));
    equaln #(12) e3589(.a(buffered_input), .b(12'b111000000101), .eq(weq3589));
    equaln #(12) e3590(.a(buffered_input), .b(12'b111000000110), .eq(weq3590));
    equaln #(12) e3591(.a(buffered_input), .b(12'b111000000111), .eq(weq3591));
    equaln #(12) e3592(.a(buffered_input), .b(12'b111000001000), .eq(weq3592));
    equaln #(12) e3593(.a(buffered_input), .b(12'b111000001001), .eq(weq3593));
    equaln #(12) e3594(.a(buffered_input), .b(12'b111000001010), .eq(weq3594));
    equaln #(12) e3595(.a(buffered_input), .b(12'b111000001011), .eq(weq3595));
    equaln #(12) e3596(.a(buffered_input), .b(12'b111000001100), .eq(weq3596));
    equaln #(12) e3597(.a(buffered_input), .b(12'b111000001101), .eq(weq3597));
    equaln #(12) e3598(.a(buffered_input), .b(12'b111000001110), .eq(weq3598));
    equaln #(12) e3599(.a(buffered_input), .b(12'b111000001111), .eq(weq3599));
    equaln #(12) e3600(.a(buffered_input), .b(12'b111000010000), .eq(weq3600));
    equaln #(12) e3601(.a(buffered_input), .b(12'b111000010001), .eq(weq3601));
    equaln #(12) e3602(.a(buffered_input), .b(12'b111000010010), .eq(weq3602));
    equaln #(12) e3603(.a(buffered_input), .b(12'b111000010011), .eq(weq3603));
    equaln #(12) e3604(.a(buffered_input), .b(12'b111000010100), .eq(weq3604));
    equaln #(12) e3605(.a(buffered_input), .b(12'b111000010101), .eq(weq3605));
    equaln #(12) e3606(.a(buffered_input), .b(12'b111000010110), .eq(weq3606));
    equaln #(12) e3607(.a(buffered_input), .b(12'b111000010111), .eq(weq3607));
    equaln #(12) e3608(.a(buffered_input), .b(12'b111000011000), .eq(weq3608));
    equaln #(12) e3609(.a(buffered_input), .b(12'b111000011001), .eq(weq3609));
    equaln #(12) e3610(.a(buffered_input), .b(12'b111000011010), .eq(weq3610));
    equaln #(12) e3611(.a(buffered_input), .b(12'b111000011011), .eq(weq3611));
    equaln #(12) e3612(.a(buffered_input), .b(12'b111000011100), .eq(weq3612));
    equaln #(12) e3613(.a(buffered_input), .b(12'b111000011101), .eq(weq3613));
    equaln #(12) e3614(.a(buffered_input), .b(12'b111000011110), .eq(weq3614));
    equaln #(12) e3615(.a(buffered_input), .b(12'b111000011111), .eq(weq3615));
    equaln #(12) e3616(.a(buffered_input), .b(12'b111000100000), .eq(weq3616));
    equaln #(12) e3617(.a(buffered_input), .b(12'b111000100001), .eq(weq3617));
    equaln #(12) e3618(.a(buffered_input), .b(12'b111000100010), .eq(weq3618));
    equaln #(12) e3619(.a(buffered_input), .b(12'b111000100011), .eq(weq3619));
    equaln #(12) e3620(.a(buffered_input), .b(12'b111000100100), .eq(weq3620));
    equaln #(12) e3621(.a(buffered_input), .b(12'b111000100101), .eq(weq3621));
    equaln #(12) e3622(.a(buffered_input), .b(12'b111000100110), .eq(weq3622));
    equaln #(12) e3623(.a(buffered_input), .b(12'b111000100111), .eq(weq3623));
    equaln #(12) e3624(.a(buffered_input), .b(12'b111000101000), .eq(weq3624));
    equaln #(12) e3625(.a(buffered_input), .b(12'b111000101001), .eq(weq3625));
    equaln #(12) e3626(.a(buffered_input), .b(12'b111000101010), .eq(weq3626));
    equaln #(12) e3627(.a(buffered_input), .b(12'b111000101011), .eq(weq3627));
    equaln #(12) e3628(.a(buffered_input), .b(12'b111000101100), .eq(weq3628));
    equaln #(12) e3629(.a(buffered_input), .b(12'b111000101101), .eq(weq3629));
    equaln #(12) e3630(.a(buffered_input), .b(12'b111000101110), .eq(weq3630));
    equaln #(12) e3631(.a(buffered_input), .b(12'b111000101111), .eq(weq3631));
    equaln #(12) e3632(.a(buffered_input), .b(12'b111000110000), .eq(weq3632));
    equaln #(12) e3633(.a(buffered_input), .b(12'b111000110001), .eq(weq3633));
    equaln #(12) e3634(.a(buffered_input), .b(12'b111000110010), .eq(weq3634));
    equaln #(12) e3635(.a(buffered_input), .b(12'b111000110011), .eq(weq3635));
    equaln #(12) e3636(.a(buffered_input), .b(12'b111000110100), .eq(weq3636));
    equaln #(12) e3637(.a(buffered_input), .b(12'b111000110101), .eq(weq3637));
    equaln #(12) e3638(.a(buffered_input), .b(12'b111000110110), .eq(weq3638));
    equaln #(12) e3639(.a(buffered_input), .b(12'b111000110111), .eq(weq3639));
    equaln #(12) e3640(.a(buffered_input), .b(12'b111000111000), .eq(weq3640));
    equaln #(12) e3641(.a(buffered_input), .b(12'b111000111001), .eq(weq3641));
    equaln #(12) e3642(.a(buffered_input), .b(12'b111000111010), .eq(weq3642));
    equaln #(12) e3643(.a(buffered_input), .b(12'b111000111011), .eq(weq3643));
    equaln #(12) e3644(.a(buffered_input), .b(12'b111000111100), .eq(weq3644));
    equaln #(12) e3645(.a(buffered_input), .b(12'b111000111101), .eq(weq3645));
    equaln #(12) e3646(.a(buffered_input), .b(12'b111000111110), .eq(weq3646));
    equaln #(12) e3647(.a(buffered_input), .b(12'b111000111111), .eq(weq3647));
    equaln #(12) e3648(.a(buffered_input), .b(12'b111001000000), .eq(weq3648));
    equaln #(12) e3649(.a(buffered_input), .b(12'b111001000001), .eq(weq3649));
    equaln #(12) e3650(.a(buffered_input), .b(12'b111001000010), .eq(weq3650));
    equaln #(12) e3651(.a(buffered_input), .b(12'b111001000011), .eq(weq3651));
    equaln #(12) e3652(.a(buffered_input), .b(12'b111001000100), .eq(weq3652));
    equaln #(12) e3653(.a(buffered_input), .b(12'b111001000101), .eq(weq3653));
    equaln #(12) e3654(.a(buffered_input), .b(12'b111001000110), .eq(weq3654));
    equaln #(12) e3655(.a(buffered_input), .b(12'b111001000111), .eq(weq3655));
    equaln #(12) e3656(.a(buffered_input), .b(12'b111001001000), .eq(weq3656));
    equaln #(12) e3657(.a(buffered_input), .b(12'b111001001001), .eq(weq3657));
    equaln #(12) e3658(.a(buffered_input), .b(12'b111001001010), .eq(weq3658));
    equaln #(12) e3659(.a(buffered_input), .b(12'b111001001011), .eq(weq3659));
    equaln #(12) e3660(.a(buffered_input), .b(12'b111001001100), .eq(weq3660));
    equaln #(12) e3661(.a(buffered_input), .b(12'b111001001101), .eq(weq3661));
    equaln #(12) e3662(.a(buffered_input), .b(12'b111001001110), .eq(weq3662));
    equaln #(12) e3663(.a(buffered_input), .b(12'b111001001111), .eq(weq3663));
    equaln #(12) e3664(.a(buffered_input), .b(12'b111001010000), .eq(weq3664));
    equaln #(12) e3665(.a(buffered_input), .b(12'b111001010001), .eq(weq3665));
    equaln #(12) e3666(.a(buffered_input), .b(12'b111001010010), .eq(weq3666));
    equaln #(12) e3667(.a(buffered_input), .b(12'b111001010011), .eq(weq3667));
    equaln #(12) e3668(.a(buffered_input), .b(12'b111001010100), .eq(weq3668));
    equaln #(12) e3669(.a(buffered_input), .b(12'b111001010101), .eq(weq3669));
    equaln #(12) e3670(.a(buffered_input), .b(12'b111001010110), .eq(weq3670));
    equaln #(12) e3671(.a(buffered_input), .b(12'b111001010111), .eq(weq3671));
    equaln #(12) e3672(.a(buffered_input), .b(12'b111001011000), .eq(weq3672));
    equaln #(12) e3673(.a(buffered_input), .b(12'b111001011001), .eq(weq3673));
    equaln #(12) e3674(.a(buffered_input), .b(12'b111001011010), .eq(weq3674));
    equaln #(12) e3675(.a(buffered_input), .b(12'b111001011011), .eq(weq3675));
    equaln #(12) e3676(.a(buffered_input), .b(12'b111001011100), .eq(weq3676));
    equaln #(12) e3677(.a(buffered_input), .b(12'b111001011101), .eq(weq3677));
    equaln #(12) e3678(.a(buffered_input), .b(12'b111001011110), .eq(weq3678));
    equaln #(12) e3679(.a(buffered_input), .b(12'b111001011111), .eq(weq3679));
    equaln #(12) e3680(.a(buffered_input), .b(12'b111001100000), .eq(weq3680));
    equaln #(12) e3681(.a(buffered_input), .b(12'b111001100001), .eq(weq3681));
    equaln #(12) e3682(.a(buffered_input), .b(12'b111001100010), .eq(weq3682));
    equaln #(12) e3683(.a(buffered_input), .b(12'b111001100011), .eq(weq3683));
    equaln #(12) e3684(.a(buffered_input), .b(12'b111001100100), .eq(weq3684));
    equaln #(12) e3685(.a(buffered_input), .b(12'b111001100101), .eq(weq3685));
    equaln #(12) e3686(.a(buffered_input), .b(12'b111001100110), .eq(weq3686));
    equaln #(12) e3687(.a(buffered_input), .b(12'b111001100111), .eq(weq3687));
    equaln #(12) e3688(.a(buffered_input), .b(12'b111001101000), .eq(weq3688));
    equaln #(12) e3689(.a(buffered_input), .b(12'b111001101001), .eq(weq3689));
    equaln #(12) e3690(.a(buffered_input), .b(12'b111001101010), .eq(weq3690));
    equaln #(12) e3691(.a(buffered_input), .b(12'b111001101011), .eq(weq3691));
    equaln #(12) e3692(.a(buffered_input), .b(12'b111001101100), .eq(weq3692));
    equaln #(12) e3693(.a(buffered_input), .b(12'b111001101101), .eq(weq3693));
    equaln #(12) e3694(.a(buffered_input), .b(12'b111001101110), .eq(weq3694));
    equaln #(12) e3695(.a(buffered_input), .b(12'b111001101111), .eq(weq3695));
    equaln #(12) e3696(.a(buffered_input), .b(12'b111001110000), .eq(weq3696));
    equaln #(12) e3697(.a(buffered_input), .b(12'b111001110001), .eq(weq3697));
    equaln #(12) e3698(.a(buffered_input), .b(12'b111001110010), .eq(weq3698));
    equaln #(12) e3699(.a(buffered_input), .b(12'b111001110011), .eq(weq3699));
    equaln #(12) e3700(.a(buffered_input), .b(12'b111001110100), .eq(weq3700));
    equaln #(12) e3701(.a(buffered_input), .b(12'b111001110101), .eq(weq3701));
    equaln #(12) e3702(.a(buffered_input), .b(12'b111001110110), .eq(weq3702));
    equaln #(12) e3703(.a(buffered_input), .b(12'b111001110111), .eq(weq3703));
    equaln #(12) e3704(.a(buffered_input), .b(12'b111001111000), .eq(weq3704));
    equaln #(12) e3705(.a(buffered_input), .b(12'b111001111001), .eq(weq3705));
    equaln #(12) e3706(.a(buffered_input), .b(12'b111001111010), .eq(weq3706));
    equaln #(12) e3707(.a(buffered_input), .b(12'b111001111011), .eq(weq3707));
    equaln #(12) e3708(.a(buffered_input), .b(12'b111001111100), .eq(weq3708));
    equaln #(12) e3709(.a(buffered_input), .b(12'b111001111101), .eq(weq3709));
    equaln #(12) e3710(.a(buffered_input), .b(12'b111001111110), .eq(weq3710));
    equaln #(12) e3711(.a(buffered_input), .b(12'b111001111111), .eq(weq3711));
    equaln #(12) e3712(.a(buffered_input), .b(12'b111010000000), .eq(weq3712));
    equaln #(12) e3713(.a(buffered_input), .b(12'b111010000001), .eq(weq3713));
    equaln #(12) e3714(.a(buffered_input), .b(12'b111010000010), .eq(weq3714));
    equaln #(12) e3715(.a(buffered_input), .b(12'b111010000011), .eq(weq3715));
    equaln #(12) e3716(.a(buffered_input), .b(12'b111010000100), .eq(weq3716));
    equaln #(12) e3717(.a(buffered_input), .b(12'b111010000101), .eq(weq3717));
    equaln #(12) e3718(.a(buffered_input), .b(12'b111010000110), .eq(weq3718));
    equaln #(12) e3719(.a(buffered_input), .b(12'b111010000111), .eq(weq3719));
    equaln #(12) e3720(.a(buffered_input), .b(12'b111010001000), .eq(weq3720));
    equaln #(12) e3721(.a(buffered_input), .b(12'b111010001001), .eq(weq3721));
    equaln #(12) e3722(.a(buffered_input), .b(12'b111010001010), .eq(weq3722));
    equaln #(12) e3723(.a(buffered_input), .b(12'b111010001011), .eq(weq3723));
    equaln #(12) e3724(.a(buffered_input), .b(12'b111010001100), .eq(weq3724));
    equaln #(12) e3725(.a(buffered_input), .b(12'b111010001101), .eq(weq3725));
    equaln #(12) e3726(.a(buffered_input), .b(12'b111010001110), .eq(weq3726));
    equaln #(12) e3727(.a(buffered_input), .b(12'b111010001111), .eq(weq3727));
    equaln #(12) e3728(.a(buffered_input), .b(12'b111010010000), .eq(weq3728));
    equaln #(12) e3729(.a(buffered_input), .b(12'b111010010001), .eq(weq3729));
    equaln #(12) e3730(.a(buffered_input), .b(12'b111010010010), .eq(weq3730));
    equaln #(12) e3731(.a(buffered_input), .b(12'b111010010011), .eq(weq3731));
    equaln #(12) e3732(.a(buffered_input), .b(12'b111010010100), .eq(weq3732));
    equaln #(12) e3733(.a(buffered_input), .b(12'b111010010101), .eq(weq3733));
    equaln #(12) e3734(.a(buffered_input), .b(12'b111010010110), .eq(weq3734));
    equaln #(12) e3735(.a(buffered_input), .b(12'b111010010111), .eq(weq3735));
    equaln #(12) e3736(.a(buffered_input), .b(12'b111010011000), .eq(weq3736));
    equaln #(12) e3737(.a(buffered_input), .b(12'b111010011001), .eq(weq3737));
    equaln #(12) e3738(.a(buffered_input), .b(12'b111010011010), .eq(weq3738));
    equaln #(12) e3739(.a(buffered_input), .b(12'b111010011011), .eq(weq3739));
    equaln #(12) e3740(.a(buffered_input), .b(12'b111010011100), .eq(weq3740));
    equaln #(12) e3741(.a(buffered_input), .b(12'b111010011101), .eq(weq3741));
    equaln #(12) e3742(.a(buffered_input), .b(12'b111010011110), .eq(weq3742));
    equaln #(12) e3743(.a(buffered_input), .b(12'b111010011111), .eq(weq3743));
    equaln #(12) e3744(.a(buffered_input), .b(12'b111010100000), .eq(weq3744));
    equaln #(12) e3745(.a(buffered_input), .b(12'b111010100001), .eq(weq3745));
    equaln #(12) e3746(.a(buffered_input), .b(12'b111010100010), .eq(weq3746));
    equaln #(12) e3747(.a(buffered_input), .b(12'b111010100011), .eq(weq3747));
    equaln #(12) e3748(.a(buffered_input), .b(12'b111010100100), .eq(weq3748));
    equaln #(12) e3749(.a(buffered_input), .b(12'b111010100101), .eq(weq3749));
    equaln #(12) e3750(.a(buffered_input), .b(12'b111010100110), .eq(weq3750));
    equaln #(12) e3751(.a(buffered_input), .b(12'b111010100111), .eq(weq3751));
    equaln #(12) e3752(.a(buffered_input), .b(12'b111010101000), .eq(weq3752));
    equaln #(12) e3753(.a(buffered_input), .b(12'b111010101001), .eq(weq3753));
    equaln #(12) e3754(.a(buffered_input), .b(12'b111010101010), .eq(weq3754));
    equaln #(12) e3755(.a(buffered_input), .b(12'b111010101011), .eq(weq3755));
    equaln #(12) e3756(.a(buffered_input), .b(12'b111010101100), .eq(weq3756));
    equaln #(12) e3757(.a(buffered_input), .b(12'b111010101101), .eq(weq3757));
    equaln #(12) e3758(.a(buffered_input), .b(12'b111010101110), .eq(weq3758));
    equaln #(12) e3759(.a(buffered_input), .b(12'b111010101111), .eq(weq3759));
    equaln #(12) e3760(.a(buffered_input), .b(12'b111010110000), .eq(weq3760));
    equaln #(12) e3761(.a(buffered_input), .b(12'b111010110001), .eq(weq3761));
    equaln #(12) e3762(.a(buffered_input), .b(12'b111010110010), .eq(weq3762));
    equaln #(12) e3763(.a(buffered_input), .b(12'b111010110011), .eq(weq3763));
    equaln #(12) e3764(.a(buffered_input), .b(12'b111010110100), .eq(weq3764));
    equaln #(12) e3765(.a(buffered_input), .b(12'b111010110101), .eq(weq3765));
    equaln #(12) e3766(.a(buffered_input), .b(12'b111010110110), .eq(weq3766));
    equaln #(12) e3767(.a(buffered_input), .b(12'b111010110111), .eq(weq3767));
    equaln #(12) e3768(.a(buffered_input), .b(12'b111010111000), .eq(weq3768));
    equaln #(12) e3769(.a(buffered_input), .b(12'b111010111001), .eq(weq3769));
    equaln #(12) e3770(.a(buffered_input), .b(12'b111010111010), .eq(weq3770));
    equaln #(12) e3771(.a(buffered_input), .b(12'b111010111011), .eq(weq3771));
    equaln #(12) e3772(.a(buffered_input), .b(12'b111010111100), .eq(weq3772));
    equaln #(12) e3773(.a(buffered_input), .b(12'b111010111101), .eq(weq3773));
    equaln #(12) e3774(.a(buffered_input), .b(12'b111010111110), .eq(weq3774));
    equaln #(12) e3775(.a(buffered_input), .b(12'b111010111111), .eq(weq3775));
    equaln #(12) e3776(.a(buffered_input), .b(12'b111011000000), .eq(weq3776));
    equaln #(12) e3777(.a(buffered_input), .b(12'b111011000001), .eq(weq3777));
    equaln #(12) e3778(.a(buffered_input), .b(12'b111011000010), .eq(weq3778));
    equaln #(12) e3779(.a(buffered_input), .b(12'b111011000011), .eq(weq3779));
    equaln #(12) e3780(.a(buffered_input), .b(12'b111011000100), .eq(weq3780));
    equaln #(12) e3781(.a(buffered_input), .b(12'b111011000101), .eq(weq3781));
    equaln #(12) e3782(.a(buffered_input), .b(12'b111011000110), .eq(weq3782));
    equaln #(12) e3783(.a(buffered_input), .b(12'b111011000111), .eq(weq3783));
    equaln #(12) e3784(.a(buffered_input), .b(12'b111011001000), .eq(weq3784));
    equaln #(12) e3785(.a(buffered_input), .b(12'b111011001001), .eq(weq3785));
    equaln #(12) e3786(.a(buffered_input), .b(12'b111011001010), .eq(weq3786));
    equaln #(12) e3787(.a(buffered_input), .b(12'b111011001011), .eq(weq3787));
    equaln #(12) e3788(.a(buffered_input), .b(12'b111011001100), .eq(weq3788));
    equaln #(12) e3789(.a(buffered_input), .b(12'b111011001101), .eq(weq3789));
    equaln #(12) e3790(.a(buffered_input), .b(12'b111011001110), .eq(weq3790));
    equaln #(12) e3791(.a(buffered_input), .b(12'b111011001111), .eq(weq3791));
    equaln #(12) e3792(.a(buffered_input), .b(12'b111011010000), .eq(weq3792));
    equaln #(12) e3793(.a(buffered_input), .b(12'b111011010001), .eq(weq3793));
    equaln #(12) e3794(.a(buffered_input), .b(12'b111011010010), .eq(weq3794));
    equaln #(12) e3795(.a(buffered_input), .b(12'b111011010011), .eq(weq3795));
    equaln #(12) e3796(.a(buffered_input), .b(12'b111011010100), .eq(weq3796));
    equaln #(12) e3797(.a(buffered_input), .b(12'b111011010101), .eq(weq3797));
    equaln #(12) e3798(.a(buffered_input), .b(12'b111011010110), .eq(weq3798));
    equaln #(12) e3799(.a(buffered_input), .b(12'b111011010111), .eq(weq3799));
    equaln #(12) e3800(.a(buffered_input), .b(12'b111011011000), .eq(weq3800));
    equaln #(12) e3801(.a(buffered_input), .b(12'b111011011001), .eq(weq3801));
    equaln #(12) e3802(.a(buffered_input), .b(12'b111011011010), .eq(weq3802));
    equaln #(12) e3803(.a(buffered_input), .b(12'b111011011011), .eq(weq3803));
    equaln #(12) e3804(.a(buffered_input), .b(12'b111011011100), .eq(weq3804));
    equaln #(12) e3805(.a(buffered_input), .b(12'b111011011101), .eq(weq3805));
    equaln #(12) e3806(.a(buffered_input), .b(12'b111011011110), .eq(weq3806));
    equaln #(12) e3807(.a(buffered_input), .b(12'b111011011111), .eq(weq3807));
    equaln #(12) e3808(.a(buffered_input), .b(12'b111011100000), .eq(weq3808));
    equaln #(12) e3809(.a(buffered_input), .b(12'b111011100001), .eq(weq3809));
    equaln #(12) e3810(.a(buffered_input), .b(12'b111011100010), .eq(weq3810));
    equaln #(12) e3811(.a(buffered_input), .b(12'b111011100011), .eq(weq3811));
    equaln #(12) e3812(.a(buffered_input), .b(12'b111011100100), .eq(weq3812));
    equaln #(12) e3813(.a(buffered_input), .b(12'b111011100101), .eq(weq3813));
    equaln #(12) e3814(.a(buffered_input), .b(12'b111011100110), .eq(weq3814));
    equaln #(12) e3815(.a(buffered_input), .b(12'b111011100111), .eq(weq3815));
    equaln #(12) e3816(.a(buffered_input), .b(12'b111011101000), .eq(weq3816));
    equaln #(12) e3817(.a(buffered_input), .b(12'b111011101001), .eq(weq3817));
    equaln #(12) e3818(.a(buffered_input), .b(12'b111011101010), .eq(weq3818));
    equaln #(12) e3819(.a(buffered_input), .b(12'b111011101011), .eq(weq3819));
    equaln #(12) e3820(.a(buffered_input), .b(12'b111011101100), .eq(weq3820));
    equaln #(12) e3821(.a(buffered_input), .b(12'b111011101101), .eq(weq3821));
    equaln #(12) e3822(.a(buffered_input), .b(12'b111011101110), .eq(weq3822));
    equaln #(12) e3823(.a(buffered_input), .b(12'b111011101111), .eq(weq3823));
    equaln #(12) e3824(.a(buffered_input), .b(12'b111011110000), .eq(weq3824));
    equaln #(12) e3825(.a(buffered_input), .b(12'b111011110001), .eq(weq3825));
    equaln #(12) e3826(.a(buffered_input), .b(12'b111011110010), .eq(weq3826));
    equaln #(12) e3827(.a(buffered_input), .b(12'b111011110011), .eq(weq3827));
    equaln #(12) e3828(.a(buffered_input), .b(12'b111011110100), .eq(weq3828));
    equaln #(12) e3829(.a(buffered_input), .b(12'b111011110101), .eq(weq3829));
    equaln #(12) e3830(.a(buffered_input), .b(12'b111011110110), .eq(weq3830));
    equaln #(12) e3831(.a(buffered_input), .b(12'b111011110111), .eq(weq3831));
    equaln #(12) e3832(.a(buffered_input), .b(12'b111011111000), .eq(weq3832));
    equaln #(12) e3833(.a(buffered_input), .b(12'b111011111001), .eq(weq3833));
    equaln #(12) e3834(.a(buffered_input), .b(12'b111011111010), .eq(weq3834));
    equaln #(12) e3835(.a(buffered_input), .b(12'b111011111011), .eq(weq3835));
    equaln #(12) e3836(.a(buffered_input), .b(12'b111011111100), .eq(weq3836));
    equaln #(12) e3837(.a(buffered_input), .b(12'b111011111101), .eq(weq3837));
    equaln #(12) e3838(.a(buffered_input), .b(12'b111011111110), .eq(weq3838));
    equaln #(12) e3839(.a(buffered_input), .b(12'b111011111111), .eq(weq3839));
    equaln #(12) e3840(.a(buffered_input), .b(12'b111100000000), .eq(weq3840));
    equaln #(12) e3841(.a(buffered_input), .b(12'b111100000001), .eq(weq3841));
    equaln #(12) e3842(.a(buffered_input), .b(12'b111100000010), .eq(weq3842));
    equaln #(12) e3843(.a(buffered_input), .b(12'b111100000011), .eq(weq3843));
    equaln #(12) e3844(.a(buffered_input), .b(12'b111100000100), .eq(weq3844));
    equaln #(12) e3845(.a(buffered_input), .b(12'b111100000101), .eq(weq3845));
    equaln #(12) e3846(.a(buffered_input), .b(12'b111100000110), .eq(weq3846));
    equaln #(12) e3847(.a(buffered_input), .b(12'b111100000111), .eq(weq3847));
    equaln #(12) e3848(.a(buffered_input), .b(12'b111100001000), .eq(weq3848));
    equaln #(12) e3849(.a(buffered_input), .b(12'b111100001001), .eq(weq3849));
    equaln #(12) e3850(.a(buffered_input), .b(12'b111100001010), .eq(weq3850));
    equaln #(12) e3851(.a(buffered_input), .b(12'b111100001011), .eq(weq3851));
    equaln #(12) e3852(.a(buffered_input), .b(12'b111100001100), .eq(weq3852));
    equaln #(12) e3853(.a(buffered_input), .b(12'b111100001101), .eq(weq3853));
    equaln #(12) e3854(.a(buffered_input), .b(12'b111100001110), .eq(weq3854));
    equaln #(12) e3855(.a(buffered_input), .b(12'b111100001111), .eq(weq3855));
    equaln #(12) e3856(.a(buffered_input), .b(12'b111100010000), .eq(weq3856));
    equaln #(12) e3857(.a(buffered_input), .b(12'b111100010001), .eq(weq3857));
    equaln #(12) e3858(.a(buffered_input), .b(12'b111100010010), .eq(weq3858));
    equaln #(12) e3859(.a(buffered_input), .b(12'b111100010011), .eq(weq3859));
    equaln #(12) e3860(.a(buffered_input), .b(12'b111100010100), .eq(weq3860));
    equaln #(12) e3861(.a(buffered_input), .b(12'b111100010101), .eq(weq3861));
    equaln #(12) e3862(.a(buffered_input), .b(12'b111100010110), .eq(weq3862));
    equaln #(12) e3863(.a(buffered_input), .b(12'b111100010111), .eq(weq3863));
    equaln #(12) e3864(.a(buffered_input), .b(12'b111100011000), .eq(weq3864));
    equaln #(12) e3865(.a(buffered_input), .b(12'b111100011001), .eq(weq3865));
    equaln #(12) e3866(.a(buffered_input), .b(12'b111100011010), .eq(weq3866));
    equaln #(12) e3867(.a(buffered_input), .b(12'b111100011011), .eq(weq3867));
    equaln #(12) e3868(.a(buffered_input), .b(12'b111100011100), .eq(weq3868));
    equaln #(12) e3869(.a(buffered_input), .b(12'b111100011101), .eq(weq3869));
    equaln #(12) e3870(.a(buffered_input), .b(12'b111100011110), .eq(weq3870));
    equaln #(12) e3871(.a(buffered_input), .b(12'b111100011111), .eq(weq3871));
    equaln #(12) e3872(.a(buffered_input), .b(12'b111100100000), .eq(weq3872));
    equaln #(12) e3873(.a(buffered_input), .b(12'b111100100001), .eq(weq3873));
    equaln #(12) e3874(.a(buffered_input), .b(12'b111100100010), .eq(weq3874));
    equaln #(12) e3875(.a(buffered_input), .b(12'b111100100011), .eq(weq3875));
    equaln #(12) e3876(.a(buffered_input), .b(12'b111100100100), .eq(weq3876));
    equaln #(12) e3877(.a(buffered_input), .b(12'b111100100101), .eq(weq3877));
    equaln #(12) e3878(.a(buffered_input), .b(12'b111100100110), .eq(weq3878));
    equaln #(12) e3879(.a(buffered_input), .b(12'b111100100111), .eq(weq3879));
    equaln #(12) e3880(.a(buffered_input), .b(12'b111100101000), .eq(weq3880));
    equaln #(12) e3881(.a(buffered_input), .b(12'b111100101001), .eq(weq3881));
    equaln #(12) e3882(.a(buffered_input), .b(12'b111100101010), .eq(weq3882));
    equaln #(12) e3883(.a(buffered_input), .b(12'b111100101011), .eq(weq3883));
    equaln #(12) e3884(.a(buffered_input), .b(12'b111100101100), .eq(weq3884));
    equaln #(12) e3885(.a(buffered_input), .b(12'b111100101101), .eq(weq3885));
    equaln #(12) e3886(.a(buffered_input), .b(12'b111100101110), .eq(weq3886));
    equaln #(12) e3887(.a(buffered_input), .b(12'b111100101111), .eq(weq3887));
    equaln #(12) e3888(.a(buffered_input), .b(12'b111100110000), .eq(weq3888));
    equaln #(12) e3889(.a(buffered_input), .b(12'b111100110001), .eq(weq3889));
    equaln #(12) e3890(.a(buffered_input), .b(12'b111100110010), .eq(weq3890));
    equaln #(12) e3891(.a(buffered_input), .b(12'b111100110011), .eq(weq3891));
    equaln #(12) e3892(.a(buffered_input), .b(12'b111100110100), .eq(weq3892));
    equaln #(12) e3893(.a(buffered_input), .b(12'b111100110101), .eq(weq3893));
    equaln #(12) e3894(.a(buffered_input), .b(12'b111100110110), .eq(weq3894));
    equaln #(12) e3895(.a(buffered_input), .b(12'b111100110111), .eq(weq3895));
    equaln #(12) e3896(.a(buffered_input), .b(12'b111100111000), .eq(weq3896));
    equaln #(12) e3897(.a(buffered_input), .b(12'b111100111001), .eq(weq3897));
    equaln #(12) e3898(.a(buffered_input), .b(12'b111100111010), .eq(weq3898));
    equaln #(12) e3899(.a(buffered_input), .b(12'b111100111011), .eq(weq3899));
    equaln #(12) e3900(.a(buffered_input), .b(12'b111100111100), .eq(weq3900));
    equaln #(12) e3901(.a(buffered_input), .b(12'b111100111101), .eq(weq3901));
    equaln #(12) e3902(.a(buffered_input), .b(12'b111100111110), .eq(weq3902));
    equaln #(12) e3903(.a(buffered_input), .b(12'b111100111111), .eq(weq3903));
    equaln #(12) e3904(.a(buffered_input), .b(12'b111101000000), .eq(weq3904));
    equaln #(12) e3905(.a(buffered_input), .b(12'b111101000001), .eq(weq3905));
    equaln #(12) e3906(.a(buffered_input), .b(12'b111101000010), .eq(weq3906));
    equaln #(12) e3907(.a(buffered_input), .b(12'b111101000011), .eq(weq3907));
    equaln #(12) e3908(.a(buffered_input), .b(12'b111101000100), .eq(weq3908));
    equaln #(12) e3909(.a(buffered_input), .b(12'b111101000101), .eq(weq3909));
    equaln #(12) e3910(.a(buffered_input), .b(12'b111101000110), .eq(weq3910));
    equaln #(12) e3911(.a(buffered_input), .b(12'b111101000111), .eq(weq3911));
    equaln #(12) e3912(.a(buffered_input), .b(12'b111101001000), .eq(weq3912));
    equaln #(12) e3913(.a(buffered_input), .b(12'b111101001001), .eq(weq3913));
    equaln #(12) e3914(.a(buffered_input), .b(12'b111101001010), .eq(weq3914));
    equaln #(12) e3915(.a(buffered_input), .b(12'b111101001011), .eq(weq3915));
    equaln #(12) e3916(.a(buffered_input), .b(12'b111101001100), .eq(weq3916));
    equaln #(12) e3917(.a(buffered_input), .b(12'b111101001101), .eq(weq3917));
    equaln #(12) e3918(.a(buffered_input), .b(12'b111101001110), .eq(weq3918));
    equaln #(12) e3919(.a(buffered_input), .b(12'b111101001111), .eq(weq3919));
    equaln #(12) e3920(.a(buffered_input), .b(12'b111101010000), .eq(weq3920));
    equaln #(12) e3921(.a(buffered_input), .b(12'b111101010001), .eq(weq3921));
    equaln #(12) e3922(.a(buffered_input), .b(12'b111101010010), .eq(weq3922));
    equaln #(12) e3923(.a(buffered_input), .b(12'b111101010011), .eq(weq3923));
    equaln #(12) e3924(.a(buffered_input), .b(12'b111101010100), .eq(weq3924));
    equaln #(12) e3925(.a(buffered_input), .b(12'b111101010101), .eq(weq3925));
    equaln #(12) e3926(.a(buffered_input), .b(12'b111101010110), .eq(weq3926));
    equaln #(12) e3927(.a(buffered_input), .b(12'b111101010111), .eq(weq3927));
    equaln #(12) e3928(.a(buffered_input), .b(12'b111101011000), .eq(weq3928));
    equaln #(12) e3929(.a(buffered_input), .b(12'b111101011001), .eq(weq3929));
    equaln #(12) e3930(.a(buffered_input), .b(12'b111101011010), .eq(weq3930));
    equaln #(12) e3931(.a(buffered_input), .b(12'b111101011011), .eq(weq3931));
    equaln #(12) e3932(.a(buffered_input), .b(12'b111101011100), .eq(weq3932));
    equaln #(12) e3933(.a(buffered_input), .b(12'b111101011101), .eq(weq3933));
    equaln #(12) e3934(.a(buffered_input), .b(12'b111101011110), .eq(weq3934));
    equaln #(12) e3935(.a(buffered_input), .b(12'b111101011111), .eq(weq3935));
    equaln #(12) e3936(.a(buffered_input), .b(12'b111101100000), .eq(weq3936));
    equaln #(12) e3937(.a(buffered_input), .b(12'b111101100001), .eq(weq3937));
    equaln #(12) e3938(.a(buffered_input), .b(12'b111101100010), .eq(weq3938));
    equaln #(12) e3939(.a(buffered_input), .b(12'b111101100011), .eq(weq3939));
    equaln #(12) e3940(.a(buffered_input), .b(12'b111101100100), .eq(weq3940));
    equaln #(12) e3941(.a(buffered_input), .b(12'b111101100101), .eq(weq3941));
    equaln #(12) e3942(.a(buffered_input), .b(12'b111101100110), .eq(weq3942));
    equaln #(12) e3943(.a(buffered_input), .b(12'b111101100111), .eq(weq3943));
    equaln #(12) e3944(.a(buffered_input), .b(12'b111101101000), .eq(weq3944));
    equaln #(12) e3945(.a(buffered_input), .b(12'b111101101001), .eq(weq3945));
    equaln #(12) e3946(.a(buffered_input), .b(12'b111101101010), .eq(weq3946));
    equaln #(12) e3947(.a(buffered_input), .b(12'b111101101011), .eq(weq3947));
    equaln #(12) e3948(.a(buffered_input), .b(12'b111101101100), .eq(weq3948));
    equaln #(12) e3949(.a(buffered_input), .b(12'b111101101101), .eq(weq3949));
    equaln #(12) e3950(.a(buffered_input), .b(12'b111101101110), .eq(weq3950));
    equaln #(12) e3951(.a(buffered_input), .b(12'b111101101111), .eq(weq3951));
    equaln #(12) e3952(.a(buffered_input), .b(12'b111101110000), .eq(weq3952));
    equaln #(12) e3953(.a(buffered_input), .b(12'b111101110001), .eq(weq3953));
    equaln #(12) e3954(.a(buffered_input), .b(12'b111101110010), .eq(weq3954));
    equaln #(12) e3955(.a(buffered_input), .b(12'b111101110011), .eq(weq3955));
    equaln #(12) e3956(.a(buffered_input), .b(12'b111101110100), .eq(weq3956));
    equaln #(12) e3957(.a(buffered_input), .b(12'b111101110101), .eq(weq3957));
    equaln #(12) e3958(.a(buffered_input), .b(12'b111101110110), .eq(weq3958));
    equaln #(12) e3959(.a(buffered_input), .b(12'b111101110111), .eq(weq3959));
    equaln #(12) e3960(.a(buffered_input), .b(12'b111101111000), .eq(weq3960));
    equaln #(12) e3961(.a(buffered_input), .b(12'b111101111001), .eq(weq3961));
    equaln #(12) e3962(.a(buffered_input), .b(12'b111101111010), .eq(weq3962));
    equaln #(12) e3963(.a(buffered_input), .b(12'b111101111011), .eq(weq3963));
    equaln #(12) e3964(.a(buffered_input), .b(12'b111101111100), .eq(weq3964));
    equaln #(12) e3965(.a(buffered_input), .b(12'b111101111101), .eq(weq3965));
    equaln #(12) e3966(.a(buffered_input), .b(12'b111101111110), .eq(weq3966));
    equaln #(12) e3967(.a(buffered_input), .b(12'b111101111111), .eq(weq3967));
    equaln #(12) e3968(.a(buffered_input), .b(12'b111110000000), .eq(weq3968));
    equaln #(12) e3969(.a(buffered_input), .b(12'b111110000001), .eq(weq3969));
    equaln #(12) e3970(.a(buffered_input), .b(12'b111110000010), .eq(weq3970));
    equaln #(12) e3971(.a(buffered_input), .b(12'b111110000011), .eq(weq3971));
    equaln #(12) e3972(.a(buffered_input), .b(12'b111110000100), .eq(weq3972));
    equaln #(12) e3973(.a(buffered_input), .b(12'b111110000101), .eq(weq3973));
    equaln #(12) e3974(.a(buffered_input), .b(12'b111110000110), .eq(weq3974));
    equaln #(12) e3975(.a(buffered_input), .b(12'b111110000111), .eq(weq3975));
    equaln #(12) e3976(.a(buffered_input), .b(12'b111110001000), .eq(weq3976));
    equaln #(12) e3977(.a(buffered_input), .b(12'b111110001001), .eq(weq3977));
    equaln #(12) e3978(.a(buffered_input), .b(12'b111110001010), .eq(weq3978));
    equaln #(12) e3979(.a(buffered_input), .b(12'b111110001011), .eq(weq3979));
    equaln #(12) e3980(.a(buffered_input), .b(12'b111110001100), .eq(weq3980));
    equaln #(12) e3981(.a(buffered_input), .b(12'b111110001101), .eq(weq3981));
    equaln #(12) e3982(.a(buffered_input), .b(12'b111110001110), .eq(weq3982));
    equaln #(12) e3983(.a(buffered_input), .b(12'b111110001111), .eq(weq3983));
    equaln #(12) e3984(.a(buffered_input), .b(12'b111110010000), .eq(weq3984));
    equaln #(12) e3985(.a(buffered_input), .b(12'b111110010001), .eq(weq3985));
    equaln #(12) e3986(.a(buffered_input), .b(12'b111110010010), .eq(weq3986));
    equaln #(12) e3987(.a(buffered_input), .b(12'b111110010011), .eq(weq3987));
    equaln #(12) e3988(.a(buffered_input), .b(12'b111110010100), .eq(weq3988));
    equaln #(12) e3989(.a(buffered_input), .b(12'b111110010101), .eq(weq3989));
    equaln #(12) e3990(.a(buffered_input), .b(12'b111110010110), .eq(weq3990));
    equaln #(12) e3991(.a(buffered_input), .b(12'b111110010111), .eq(weq3991));
    equaln #(12) e3992(.a(buffered_input), .b(12'b111110011000), .eq(weq3992));
    equaln #(12) e3993(.a(buffered_input), .b(12'b111110011001), .eq(weq3993));
    equaln #(12) e3994(.a(buffered_input), .b(12'b111110011010), .eq(weq3994));
    equaln #(12) e3995(.a(buffered_input), .b(12'b111110011011), .eq(weq3995));
    equaln #(12) e3996(.a(buffered_input), .b(12'b111110011100), .eq(weq3996));
    equaln #(12) e3997(.a(buffered_input), .b(12'b111110011101), .eq(weq3997));
    equaln #(12) e3998(.a(buffered_input), .b(12'b111110011110), .eq(weq3998));
    equaln #(12) e3999(.a(buffered_input), .b(12'b111110011111), .eq(weq3999));
    equaln #(12) e4000(.a(buffered_input), .b(12'b111110100000), .eq(weq4000));
    equaln #(12) e4001(.a(buffered_input), .b(12'b111110100001), .eq(weq4001));
    equaln #(12) e4002(.a(buffered_input), .b(12'b111110100010), .eq(weq4002));
    equaln #(12) e4003(.a(buffered_input), .b(12'b111110100011), .eq(weq4003));
    equaln #(12) e4004(.a(buffered_input), .b(12'b111110100100), .eq(weq4004));
    equaln #(12) e4005(.a(buffered_input), .b(12'b111110100101), .eq(weq4005));
    equaln #(12) e4006(.a(buffered_input), .b(12'b111110100110), .eq(weq4006));
    equaln #(12) e4007(.a(buffered_input), .b(12'b111110100111), .eq(weq4007));
    equaln #(12) e4008(.a(buffered_input), .b(12'b111110101000), .eq(weq4008));
    equaln #(12) e4009(.a(buffered_input), .b(12'b111110101001), .eq(weq4009));
    equaln #(12) e4010(.a(buffered_input), .b(12'b111110101010), .eq(weq4010));
    equaln #(12) e4011(.a(buffered_input), .b(12'b111110101011), .eq(weq4011));
    equaln #(12) e4012(.a(buffered_input), .b(12'b111110101100), .eq(weq4012));
    equaln #(12) e4013(.a(buffered_input), .b(12'b111110101101), .eq(weq4013));
    equaln #(12) e4014(.a(buffered_input), .b(12'b111110101110), .eq(weq4014));
    equaln #(12) e4015(.a(buffered_input), .b(12'b111110101111), .eq(weq4015));
    equaln #(12) e4016(.a(buffered_input), .b(12'b111110110000), .eq(weq4016));
    equaln #(12) e4017(.a(buffered_input), .b(12'b111110110001), .eq(weq4017));
    equaln #(12) e4018(.a(buffered_input), .b(12'b111110110010), .eq(weq4018));
    equaln #(12) e4019(.a(buffered_input), .b(12'b111110110011), .eq(weq4019));
    equaln #(12) e4020(.a(buffered_input), .b(12'b111110110100), .eq(weq4020));
    equaln #(12) e4021(.a(buffered_input), .b(12'b111110110101), .eq(weq4021));
    equaln #(12) e4022(.a(buffered_input), .b(12'b111110110110), .eq(weq4022));
    equaln #(12) e4023(.a(buffered_input), .b(12'b111110110111), .eq(weq4023));
    equaln #(12) e4024(.a(buffered_input), .b(12'b111110111000), .eq(weq4024));
    equaln #(12) e4025(.a(buffered_input), .b(12'b111110111001), .eq(weq4025));
    equaln #(12) e4026(.a(buffered_input), .b(12'b111110111010), .eq(weq4026));
    equaln #(12) e4027(.a(buffered_input), .b(12'b111110111011), .eq(weq4027));
    equaln #(12) e4028(.a(buffered_input), .b(12'b111110111100), .eq(weq4028));
    equaln #(12) e4029(.a(buffered_input), .b(12'b111110111101), .eq(weq4029));
    equaln #(12) e4030(.a(buffered_input), .b(12'b111110111110), .eq(weq4030));
    equaln #(12) e4031(.a(buffered_input), .b(12'b111110111111), .eq(weq4031));
    equaln #(12) e4032(.a(buffered_input), .b(12'b111111000000), .eq(weq4032));
    equaln #(12) e4033(.a(buffered_input), .b(12'b111111000001), .eq(weq4033));
    equaln #(12) e4034(.a(buffered_input), .b(12'b111111000010), .eq(weq4034));
    equaln #(12) e4035(.a(buffered_input), .b(12'b111111000011), .eq(weq4035));
    equaln #(12) e4036(.a(buffered_input), .b(12'b111111000100), .eq(weq4036));
    equaln #(12) e4037(.a(buffered_input), .b(12'b111111000101), .eq(weq4037));
    equaln #(12) e4038(.a(buffered_input), .b(12'b111111000110), .eq(weq4038));
    equaln #(12) e4039(.a(buffered_input), .b(12'b111111000111), .eq(weq4039));
    equaln #(12) e4040(.a(buffered_input), .b(12'b111111001000), .eq(weq4040));
    equaln #(12) e4041(.a(buffered_input), .b(12'b111111001001), .eq(weq4041));
    equaln #(12) e4042(.a(buffered_input), .b(12'b111111001010), .eq(weq4042));
    equaln #(12) e4043(.a(buffered_input), .b(12'b111111001011), .eq(weq4043));
    equaln #(12) e4044(.a(buffered_input), .b(12'b111111001100), .eq(weq4044));
    equaln #(12) e4045(.a(buffered_input), .b(12'b111111001101), .eq(weq4045));
    equaln #(12) e4046(.a(buffered_input), .b(12'b111111001110), .eq(weq4046));
    equaln #(12) e4047(.a(buffered_input), .b(12'b111111001111), .eq(weq4047));
    equaln #(12) e4048(.a(buffered_input), .b(12'b111111010000), .eq(weq4048));
    equaln #(12) e4049(.a(buffered_input), .b(12'b111111010001), .eq(weq4049));
    equaln #(12) e4050(.a(buffered_input), .b(12'b111111010010), .eq(weq4050));
    equaln #(12) e4051(.a(buffered_input), .b(12'b111111010011), .eq(weq4051));
    equaln #(12) e4052(.a(buffered_input), .b(12'b111111010100), .eq(weq4052));
    equaln #(12) e4053(.a(buffered_input), .b(12'b111111010101), .eq(weq4053));
    equaln #(12) e4054(.a(buffered_input), .b(12'b111111010110), .eq(weq4054));
    equaln #(12) e4055(.a(buffered_input), .b(12'b111111010111), .eq(weq4055));
    equaln #(12) e4056(.a(buffered_input), .b(12'b111111011000), .eq(weq4056));
    equaln #(12) e4057(.a(buffered_input), .b(12'b111111011001), .eq(weq4057));
    equaln #(12) e4058(.a(buffered_input), .b(12'b111111011010), .eq(weq4058));
    equaln #(12) e4059(.a(buffered_input), .b(12'b111111011011), .eq(weq4059));
    equaln #(12) e4060(.a(buffered_input), .b(12'b111111011100), .eq(weq4060));
    equaln #(12) e4061(.a(buffered_input), .b(12'b111111011101), .eq(weq4061));
    equaln #(12) e4062(.a(buffered_input), .b(12'b111111011110), .eq(weq4062));
    equaln #(12) e4063(.a(buffered_input), .b(12'b111111011111), .eq(weq4063));
    equaln #(12) e4064(.a(buffered_input), .b(12'b111111100000), .eq(weq4064));
    equaln #(12) e4065(.a(buffered_input), .b(12'b111111100001), .eq(weq4065));
    equaln #(12) e4066(.a(buffered_input), .b(12'b111111100010), .eq(weq4066));
    equaln #(12) e4067(.a(buffered_input), .b(12'b111111100011), .eq(weq4067));
    equaln #(12) e4068(.a(buffered_input), .b(12'b111111100100), .eq(weq4068));
    equaln #(12) e4069(.a(buffered_input), .b(12'b111111100101), .eq(weq4069));
    equaln #(12) e4070(.a(buffered_input), .b(12'b111111100110), .eq(weq4070));
    equaln #(12) e4071(.a(buffered_input), .b(12'b111111100111), .eq(weq4071));
    equaln #(12) e4072(.a(buffered_input), .b(12'b111111101000), .eq(weq4072));
    equaln #(12) e4073(.a(buffered_input), .b(12'b111111101001), .eq(weq4073));
    equaln #(12) e4074(.a(buffered_input), .b(12'b111111101010), .eq(weq4074));
    equaln #(12) e4075(.a(buffered_input), .b(12'b111111101011), .eq(weq4075));
    equaln #(12) e4076(.a(buffered_input), .b(12'b111111101100), .eq(weq4076));
    equaln #(12) e4077(.a(buffered_input), .b(12'b111111101101), .eq(weq4077));
    equaln #(12) e4078(.a(buffered_input), .b(12'b111111101110), .eq(weq4078));
    equaln #(12) e4079(.a(buffered_input), .b(12'b111111101111), .eq(weq4079));
    equaln #(12) e4080(.a(buffered_input), .b(12'b111111110000), .eq(weq4080));
    equaln #(12) e4081(.a(buffered_input), .b(12'b111111110001), .eq(weq4081));
    equaln #(12) e4082(.a(buffered_input), .b(12'b111111110010), .eq(weq4082));
    equaln #(12) e4083(.a(buffered_input), .b(12'b111111110011), .eq(weq4083));
    equaln #(12) e4084(.a(buffered_input), .b(12'b111111110100), .eq(weq4084));
    equaln #(12) e4085(.a(buffered_input), .b(12'b111111110101), .eq(weq4085));
    equaln #(12) e4086(.a(buffered_input), .b(12'b111111110110), .eq(weq4086));
    equaln #(12) e4087(.a(buffered_input), .b(12'b111111110111), .eq(weq4087));
    equaln #(12) e4088(.a(buffered_input), .b(12'b111111111000), .eq(weq4088));
    equaln #(12) e4089(.a(buffered_input), .b(12'b111111111001), .eq(weq4089));
    equaln #(12) e4090(.a(buffered_input), .b(12'b111111111010), .eq(weq4090));
    equaln #(12) e4091(.a(buffered_input), .b(12'b111111111011), .eq(weq4091));
    equaln #(12) e4092(.a(buffered_input), .b(12'b111111111100), .eq(weq4092));
    equaln #(12) e4093(.a(buffered_input), .b(12'b111111111101), .eq(weq4093));
    equaln #(12) e4094(.a(buffered_input), .b(12'b111111111110), .eq(weq4094));
    equaln #(12) e4095(.a(buffered_input), .b(12'b111111111111), .eq(weq4095));
    assign out = {weq4095, weq4094, weq4093, weq4092, weq4091, weq4090, weq4089, weq4088, weq4087, weq4086, weq4085, weq4084, weq4083, weq4082, weq4081, weq4080, weq4079, weq4078, weq4077, weq4076, weq4075, weq4074, weq4073, weq4072, weq4071, weq4070, weq4069, weq4068, weq4067, weq4066, weq4065, weq4064, weq4063, weq4062, weq4061, weq4060, weq4059, weq4058, weq4057, weq4056, weq4055, weq4054, weq4053, weq4052, weq4051, weq4050, weq4049, weq4048, weq4047, weq4046, weq4045, weq4044, weq4043, weq4042, weq4041, weq4040, weq4039, weq4038, weq4037, weq4036, weq4035, weq4034, weq4033, weq4032, weq4031, weq4030, weq4029, weq4028, weq4027, weq4026, weq4025, weq4024, weq4023, weq4022, weq4021, weq4020, weq4019, weq4018, weq4017, weq4016, weq4015, weq4014, weq4013, weq4012, weq4011, weq4010, weq4009, weq4008, weq4007, weq4006, weq4005, weq4004, weq4003, weq4002, weq4001, weq4000, weq3999, weq3998, weq3997, weq3996, weq3995, weq3994, weq3993, weq3992, weq3991, weq3990, weq3989, weq3988, weq3987, weq3986, weq3985, weq3984, weq3983, weq3982, weq3981, weq3980, weq3979, weq3978, weq3977, weq3976, weq3975, weq3974, weq3973, weq3972, weq3971, weq3970, weq3969, weq3968, weq3967, weq3966, weq3965, weq3964, weq3963, weq3962, weq3961, weq3960, weq3959, weq3958, weq3957, weq3956, weq3955, weq3954, weq3953, weq3952, weq3951, weq3950, weq3949, weq3948, weq3947, weq3946, weq3945, weq3944, weq3943, weq3942, weq3941, weq3940, weq3939, weq3938, weq3937, weq3936, weq3935, weq3934, weq3933, weq3932, weq3931, weq3930, weq3929, weq3928, weq3927, weq3926, weq3925, weq3924, weq3923, weq3922, weq3921, weq3920, weq3919, weq3918, weq3917, weq3916, weq3915, weq3914, weq3913, weq3912, weq3911, weq3910, weq3909, weq3908, weq3907, weq3906, weq3905, weq3904, weq3903, weq3902, weq3901, weq3900, weq3899, weq3898, weq3897, weq3896, weq3895, weq3894, weq3893, weq3892, weq3891, weq3890, weq3889, weq3888, weq3887, weq3886, weq3885, weq3884, weq3883, weq3882, weq3881, weq3880, weq3879, weq3878, weq3877, weq3876, weq3875, weq3874, weq3873, weq3872, weq3871, weq3870, weq3869, weq3868, weq3867, weq3866, weq3865, weq3864, weq3863, weq3862, weq3861, weq3860, weq3859, weq3858, weq3857, weq3856, weq3855, weq3854, weq3853, weq3852, weq3851, weq3850, weq3849, weq3848, weq3847, weq3846, weq3845, weq3844, weq3843, weq3842, weq3841, weq3840, weq3839, weq3838, weq3837, weq3836, weq3835, weq3834, weq3833, weq3832, weq3831, weq3830, weq3829, weq3828, weq3827, weq3826, weq3825, weq3824, weq3823, weq3822, weq3821, weq3820, weq3819, weq3818, weq3817, weq3816, weq3815, weq3814, weq3813, weq3812, weq3811, weq3810, weq3809, weq3808, weq3807, weq3806, weq3805, weq3804, weq3803, weq3802, weq3801, weq3800, weq3799, weq3798, weq3797, weq3796, weq3795, weq3794, weq3793, weq3792, weq3791, weq3790, weq3789, weq3788, weq3787, weq3786, weq3785, weq3784, weq3783, weq3782, weq3781, weq3780, weq3779, weq3778, weq3777, weq3776, weq3775, weq3774, weq3773, weq3772, weq3771, weq3770, weq3769, weq3768, weq3767, weq3766, weq3765, weq3764, weq3763, weq3762, weq3761, weq3760, weq3759, weq3758, weq3757, weq3756, weq3755, weq3754, weq3753, weq3752, weq3751, weq3750, weq3749, weq3748, weq3747, weq3746, weq3745, weq3744, weq3743, weq3742, weq3741, weq3740, weq3739, weq3738, weq3737, weq3736, weq3735, weq3734, weq3733, weq3732, weq3731, weq3730, weq3729, weq3728, weq3727, weq3726, weq3725, weq3724, weq3723, weq3722, weq3721, weq3720, weq3719, weq3718, weq3717, weq3716, weq3715, weq3714, weq3713, weq3712, weq3711, weq3710, weq3709, weq3708, weq3707, weq3706, weq3705, weq3704, weq3703, weq3702, weq3701, weq3700, weq3699, weq3698, weq3697, weq3696, weq3695, weq3694, weq3693, weq3692, weq3691, weq3690, weq3689, weq3688, weq3687, weq3686, weq3685, weq3684, weq3683, weq3682, weq3681, weq3680, weq3679, weq3678, weq3677, weq3676, weq3675, weq3674, weq3673, weq3672, weq3671, weq3670, weq3669, weq3668, weq3667, weq3666, weq3665, weq3664, weq3663, weq3662, weq3661, weq3660, weq3659, weq3658, weq3657, weq3656, weq3655, weq3654, weq3653, weq3652, weq3651, weq3650, weq3649, weq3648, weq3647, weq3646, weq3645, weq3644, weq3643, weq3642, weq3641, weq3640, weq3639, weq3638, weq3637, weq3636, weq3635, weq3634, weq3633, weq3632, weq3631, weq3630, weq3629, weq3628, weq3627, weq3626, weq3625, weq3624, weq3623, weq3622, weq3621, weq3620, weq3619, weq3618, weq3617, weq3616, weq3615, weq3614, weq3613, weq3612, weq3611, weq3610, weq3609, weq3608, weq3607, weq3606, weq3605, weq3604, weq3603, weq3602, weq3601, weq3600, weq3599, weq3598, weq3597, weq3596, weq3595, weq3594, weq3593, weq3592, weq3591, weq3590, weq3589, weq3588, weq3587, weq3586, weq3585, weq3584, weq3583, weq3582, weq3581, weq3580, weq3579, weq3578, weq3577, weq3576, weq3575, weq3574, weq3573, weq3572, weq3571, weq3570, weq3569, weq3568, weq3567, weq3566, weq3565, weq3564, weq3563, weq3562, weq3561, weq3560, weq3559, weq3558, weq3557, weq3556, weq3555, weq3554, weq3553, weq3552, weq3551, weq3550, weq3549, weq3548, weq3547, weq3546, weq3545, weq3544, weq3543, weq3542, weq3541, weq3540, weq3539, weq3538, weq3537, weq3536, weq3535, weq3534, weq3533, weq3532, weq3531, weq3530, weq3529, weq3528, weq3527, weq3526, weq3525, weq3524, weq3523, weq3522, weq3521, weq3520, weq3519, weq3518, weq3517, weq3516, weq3515, weq3514, weq3513, weq3512, weq3511, weq3510, weq3509, weq3508, weq3507, weq3506, weq3505, weq3504, weq3503, weq3502, weq3501, weq3500, weq3499, weq3498, weq3497, weq3496, weq3495, weq3494, weq3493, weq3492, weq3491, weq3490, weq3489, weq3488, weq3487, weq3486, weq3485, weq3484, weq3483, weq3482, weq3481, weq3480, weq3479, weq3478, weq3477, weq3476, weq3475, weq3474, weq3473, weq3472, weq3471, weq3470, weq3469, weq3468, weq3467, weq3466, weq3465, weq3464, weq3463, weq3462, weq3461, weq3460, weq3459, weq3458, weq3457, weq3456, weq3455, weq3454, weq3453, weq3452, weq3451, weq3450, weq3449, weq3448, weq3447, weq3446, weq3445, weq3444, weq3443, weq3442, weq3441, weq3440, weq3439, weq3438, weq3437, weq3436, weq3435, weq3434, weq3433, weq3432, weq3431, weq3430, weq3429, weq3428, weq3427, weq3426, weq3425, weq3424, weq3423, weq3422, weq3421, weq3420, weq3419, weq3418, weq3417, weq3416, weq3415, weq3414, weq3413, weq3412, weq3411, weq3410, weq3409, weq3408, weq3407, weq3406, weq3405, weq3404, weq3403, weq3402, weq3401, weq3400, weq3399, weq3398, weq3397, weq3396, weq3395, weq3394, weq3393, weq3392, weq3391, weq3390, weq3389, weq3388, weq3387, weq3386, weq3385, weq3384, weq3383, weq3382, weq3381, weq3380, weq3379, weq3378, weq3377, weq3376, weq3375, weq3374, weq3373, weq3372, weq3371, weq3370, weq3369, weq3368, weq3367, weq3366, weq3365, weq3364, weq3363, weq3362, weq3361, weq3360, weq3359, weq3358, weq3357, weq3356, weq3355, weq3354, weq3353, weq3352, weq3351, weq3350, weq3349, weq3348, weq3347, weq3346, weq3345, weq3344, weq3343, weq3342, weq3341, weq3340, weq3339, weq3338, weq3337, weq3336, weq3335, weq3334, weq3333, weq3332, weq3331, weq3330, weq3329, weq3328, weq3327, weq3326, weq3325, weq3324, weq3323, weq3322, weq3321, weq3320, weq3319, weq3318, weq3317, weq3316, weq3315, weq3314, weq3313, weq3312, weq3311, weq3310, weq3309, weq3308, weq3307, weq3306, weq3305, weq3304, weq3303, weq3302, weq3301, weq3300, weq3299, weq3298, weq3297, weq3296, weq3295, weq3294, weq3293, weq3292, weq3291, weq3290, weq3289, weq3288, weq3287, weq3286, weq3285, weq3284, weq3283, weq3282, weq3281, weq3280, weq3279, weq3278, weq3277, weq3276, weq3275, weq3274, weq3273, weq3272, weq3271, weq3270, weq3269, weq3268, weq3267, weq3266, weq3265, weq3264, weq3263, weq3262, weq3261, weq3260, weq3259, weq3258, weq3257, weq3256, weq3255, weq3254, weq3253, weq3252, weq3251, weq3250, weq3249, weq3248, weq3247, weq3246, weq3245, weq3244, weq3243, weq3242, weq3241, weq3240, weq3239, weq3238, weq3237, weq3236, weq3235, weq3234, weq3233, weq3232, weq3231, weq3230, weq3229, weq3228, weq3227, weq3226, weq3225, weq3224, weq3223, weq3222, weq3221, weq3220, weq3219, weq3218, weq3217, weq3216, weq3215, weq3214, weq3213, weq3212, weq3211, weq3210, weq3209, weq3208, weq3207, weq3206, weq3205, weq3204, weq3203, weq3202, weq3201, weq3200, weq3199, weq3198, weq3197, weq3196, weq3195, weq3194, weq3193, weq3192, weq3191, weq3190, weq3189, weq3188, weq3187, weq3186, weq3185, weq3184, weq3183, weq3182, weq3181, weq3180, weq3179, weq3178, weq3177, weq3176, weq3175, weq3174, weq3173, weq3172, weq3171, weq3170, weq3169, weq3168, weq3167, weq3166, weq3165, weq3164, weq3163, weq3162, weq3161, weq3160, weq3159, weq3158, weq3157, weq3156, weq3155, weq3154, weq3153, weq3152, weq3151, weq3150, weq3149, weq3148, weq3147, weq3146, weq3145, weq3144, weq3143, weq3142, weq3141, weq3140, weq3139, weq3138, weq3137, weq3136, weq3135, weq3134, weq3133, weq3132, weq3131, weq3130, weq3129, weq3128, weq3127, weq3126, weq3125, weq3124, weq3123, weq3122, weq3121, weq3120, weq3119, weq3118, weq3117, weq3116, weq3115, weq3114, weq3113, weq3112, weq3111, weq3110, weq3109, weq3108, weq3107, weq3106, weq3105, weq3104, weq3103, weq3102, weq3101, weq3100, weq3099, weq3098, weq3097, weq3096, weq3095, weq3094, weq3093, weq3092, weq3091, weq3090, weq3089, weq3088, weq3087, weq3086, weq3085, weq3084, weq3083, weq3082, weq3081, weq3080, weq3079, weq3078, weq3077, weq3076, weq3075, weq3074, weq3073, weq3072, weq3071, weq3070, weq3069, weq3068, weq3067, weq3066, weq3065, weq3064, weq3063, weq3062, weq3061, weq3060, weq3059, weq3058, weq3057, weq3056, weq3055, weq3054, weq3053, weq3052, weq3051, weq3050, weq3049, weq3048, weq3047, weq3046, weq3045, weq3044, weq3043, weq3042, weq3041, weq3040, weq3039, weq3038, weq3037, weq3036, weq3035, weq3034, weq3033, weq3032, weq3031, weq3030, weq3029, weq3028, weq3027, weq3026, weq3025, weq3024, weq3023, weq3022, weq3021, weq3020, weq3019, weq3018, weq3017, weq3016, weq3015, weq3014, weq3013, weq3012, weq3011, weq3010, weq3009, weq3008, weq3007, weq3006, weq3005, weq3004, weq3003, weq3002, weq3001, weq3000, weq2999, weq2998, weq2997, weq2996, weq2995, weq2994, weq2993, weq2992, weq2991, weq2990, weq2989, weq2988, weq2987, weq2986, weq2985, weq2984, weq2983, weq2982, weq2981, weq2980, weq2979, weq2978, weq2977, weq2976, weq2975, weq2974, weq2973, weq2972, weq2971, weq2970, weq2969, weq2968, weq2967, weq2966, weq2965, weq2964, weq2963, weq2962, weq2961, weq2960, weq2959, weq2958, weq2957, weq2956, weq2955, weq2954, weq2953, weq2952, weq2951, weq2950, weq2949, weq2948, weq2947, weq2946, weq2945, weq2944, weq2943, weq2942, weq2941, weq2940, weq2939, weq2938, weq2937, weq2936, weq2935, weq2934, weq2933, weq2932, weq2931, weq2930, weq2929, weq2928, weq2927, weq2926, weq2925, weq2924, weq2923, weq2922, weq2921, weq2920, weq2919, weq2918, weq2917, weq2916, weq2915, weq2914, weq2913, weq2912, weq2911, weq2910, weq2909, weq2908, weq2907, weq2906, weq2905, weq2904, weq2903, weq2902, weq2901, weq2900, weq2899, weq2898, weq2897, weq2896, weq2895, weq2894, weq2893, weq2892, weq2891, weq2890, weq2889, weq2888, weq2887, weq2886, weq2885, weq2884, weq2883, weq2882, weq2881, weq2880, weq2879, weq2878, weq2877, weq2876, weq2875, weq2874, weq2873, weq2872, weq2871, weq2870, weq2869, weq2868, weq2867, weq2866, weq2865, weq2864, weq2863, weq2862, weq2861, weq2860, weq2859, weq2858, weq2857, weq2856, weq2855, weq2854, weq2853, weq2852, weq2851, weq2850, weq2849, weq2848, weq2847, weq2846, weq2845, weq2844, weq2843, weq2842, weq2841, weq2840, weq2839, weq2838, weq2837, weq2836, weq2835, weq2834, weq2833, weq2832, weq2831, weq2830, weq2829, weq2828, weq2827, weq2826, weq2825, weq2824, weq2823, weq2822, weq2821, weq2820, weq2819, weq2818, weq2817, weq2816, weq2815, weq2814, weq2813, weq2812, weq2811, weq2810, weq2809, weq2808, weq2807, weq2806, weq2805, weq2804, weq2803, weq2802, weq2801, weq2800, weq2799, weq2798, weq2797, weq2796, weq2795, weq2794, weq2793, weq2792, weq2791, weq2790, weq2789, weq2788, weq2787, weq2786, weq2785, weq2784, weq2783, weq2782, weq2781, weq2780, weq2779, weq2778, weq2777, weq2776, weq2775, weq2774, weq2773, weq2772, weq2771, weq2770, weq2769, weq2768, weq2767, weq2766, weq2765, weq2764, weq2763, weq2762, weq2761, weq2760, weq2759, weq2758, weq2757, weq2756, weq2755, weq2754, weq2753, weq2752, weq2751, weq2750, weq2749, weq2748, weq2747, weq2746, weq2745, weq2744, weq2743, weq2742, weq2741, weq2740, weq2739, weq2738, weq2737, weq2736, weq2735, weq2734, weq2733, weq2732, weq2731, weq2730, weq2729, weq2728, weq2727, weq2726, weq2725, weq2724, weq2723, weq2722, weq2721, weq2720, weq2719, weq2718, weq2717, weq2716, weq2715, weq2714, weq2713, weq2712, weq2711, weq2710, weq2709, weq2708, weq2707, weq2706, weq2705, weq2704, weq2703, weq2702, weq2701, weq2700, weq2699, weq2698, weq2697, weq2696, weq2695, weq2694, weq2693, weq2692, weq2691, weq2690, weq2689, weq2688, weq2687, weq2686, weq2685, weq2684, weq2683, weq2682, weq2681, weq2680, weq2679, weq2678, weq2677, weq2676, weq2675, weq2674, weq2673, weq2672, weq2671, weq2670, weq2669, weq2668, weq2667, weq2666, weq2665, weq2664, weq2663, weq2662, weq2661, weq2660, weq2659, weq2658, weq2657, weq2656, weq2655, weq2654, weq2653, weq2652, weq2651, weq2650, weq2649, weq2648, weq2647, weq2646, weq2645, weq2644, weq2643, weq2642, weq2641, weq2640, weq2639, weq2638, weq2637, weq2636, weq2635, weq2634, weq2633, weq2632, weq2631, weq2630, weq2629, weq2628, weq2627, weq2626, weq2625, weq2624, weq2623, weq2622, weq2621, weq2620, weq2619, weq2618, weq2617, weq2616, weq2615, weq2614, weq2613, weq2612, weq2611, weq2610, weq2609, weq2608, weq2607, weq2606, weq2605, weq2604, weq2603, weq2602, weq2601, weq2600, weq2599, weq2598, weq2597, weq2596, weq2595, weq2594, weq2593, weq2592, weq2591, weq2590, weq2589, weq2588, weq2587, weq2586, weq2585, weq2584, weq2583, weq2582, weq2581, weq2580, weq2579, weq2578, weq2577, weq2576, weq2575, weq2574, weq2573, weq2572, weq2571, weq2570, weq2569, weq2568, weq2567, weq2566, weq2565, weq2564, weq2563, weq2562, weq2561, weq2560, weq2559, weq2558, weq2557, weq2556, weq2555, weq2554, weq2553, weq2552, weq2551, weq2550, weq2549, weq2548, weq2547, weq2546, weq2545, weq2544, weq2543, weq2542, weq2541, weq2540, weq2539, weq2538, weq2537, weq2536, weq2535, weq2534, weq2533, weq2532, weq2531, weq2530, weq2529, weq2528, weq2527, weq2526, weq2525, weq2524, weq2523, weq2522, weq2521, weq2520, weq2519, weq2518, weq2517, weq2516, weq2515, weq2514, weq2513, weq2512, weq2511, weq2510, weq2509, weq2508, weq2507, weq2506, weq2505, weq2504, weq2503, weq2502, weq2501, weq2500, weq2499, weq2498, weq2497, weq2496, weq2495, weq2494, weq2493, weq2492, weq2491, weq2490, weq2489, weq2488, weq2487, weq2486, weq2485, weq2484, weq2483, weq2482, weq2481, weq2480, weq2479, weq2478, weq2477, weq2476, weq2475, weq2474, weq2473, weq2472, weq2471, weq2470, weq2469, weq2468, weq2467, weq2466, weq2465, weq2464, weq2463, weq2462, weq2461, weq2460, weq2459, weq2458, weq2457, weq2456, weq2455, weq2454, weq2453, weq2452, weq2451, weq2450, weq2449, weq2448, weq2447, weq2446, weq2445, weq2444, weq2443, weq2442, weq2441, weq2440, weq2439, weq2438, weq2437, weq2436, weq2435, weq2434, weq2433, weq2432, weq2431, weq2430, weq2429, weq2428, weq2427, weq2426, weq2425, weq2424, weq2423, weq2422, weq2421, weq2420, weq2419, weq2418, weq2417, weq2416, weq2415, weq2414, weq2413, weq2412, weq2411, weq2410, weq2409, weq2408, weq2407, weq2406, weq2405, weq2404, weq2403, weq2402, weq2401, weq2400, weq2399, weq2398, weq2397, weq2396, weq2395, weq2394, weq2393, weq2392, weq2391, weq2390, weq2389, weq2388, weq2387, weq2386, weq2385, weq2384, weq2383, weq2382, weq2381, weq2380, weq2379, weq2378, weq2377, weq2376, weq2375, weq2374, weq2373, weq2372, weq2371, weq2370, weq2369, weq2368, weq2367, weq2366, weq2365, weq2364, weq2363, weq2362, weq2361, weq2360, weq2359, weq2358, weq2357, weq2356, weq2355, weq2354, weq2353, weq2352, weq2351, weq2350, weq2349, weq2348, weq2347, weq2346, weq2345, weq2344, weq2343, weq2342, weq2341, weq2340, weq2339, weq2338, weq2337, weq2336, weq2335, weq2334, weq2333, weq2332, weq2331, weq2330, weq2329, weq2328, weq2327, weq2326, weq2325, weq2324, weq2323, weq2322, weq2321, weq2320, weq2319, weq2318, weq2317, weq2316, weq2315, weq2314, weq2313, weq2312, weq2311, weq2310, weq2309, weq2308, weq2307, weq2306, weq2305, weq2304, weq2303, weq2302, weq2301, weq2300, weq2299, weq2298, weq2297, weq2296, weq2295, weq2294, weq2293, weq2292, weq2291, weq2290, weq2289, weq2288, weq2287, weq2286, weq2285, weq2284, weq2283, weq2282, weq2281, weq2280, weq2279, weq2278, weq2277, weq2276, weq2275, weq2274, weq2273, weq2272, weq2271, weq2270, weq2269, weq2268, weq2267, weq2266, weq2265, weq2264, weq2263, weq2262, weq2261, weq2260, weq2259, weq2258, weq2257, weq2256, weq2255, weq2254, weq2253, weq2252, weq2251, weq2250, weq2249, weq2248, weq2247, weq2246, weq2245, weq2244, weq2243, weq2242, weq2241, weq2240, weq2239, weq2238, weq2237, weq2236, weq2235, weq2234, weq2233, weq2232, weq2231, weq2230, weq2229, weq2228, weq2227, weq2226, weq2225, weq2224, weq2223, weq2222, weq2221, weq2220, weq2219, weq2218, weq2217, weq2216, weq2215, weq2214, weq2213, weq2212, weq2211, weq2210, weq2209, weq2208, weq2207, weq2206, weq2205, weq2204, weq2203, weq2202, weq2201, weq2200, weq2199, weq2198, weq2197, weq2196, weq2195, weq2194, weq2193, weq2192, weq2191, weq2190, weq2189, weq2188, weq2187, weq2186, weq2185, weq2184, weq2183, weq2182, weq2181, weq2180, weq2179, weq2178, weq2177, weq2176, weq2175, weq2174, weq2173, weq2172, weq2171, weq2170, weq2169, weq2168, weq2167, weq2166, weq2165, weq2164, weq2163, weq2162, weq2161, weq2160, weq2159, weq2158, weq2157, weq2156, weq2155, weq2154, weq2153, weq2152, weq2151, weq2150, weq2149, weq2148, weq2147, weq2146, weq2145, weq2144, weq2143, weq2142, weq2141, weq2140, weq2139, weq2138, weq2137, weq2136, weq2135, weq2134, weq2133, weq2132, weq2131, weq2130, weq2129, weq2128, weq2127, weq2126, weq2125, weq2124, weq2123, weq2122, weq2121, weq2120, weq2119, weq2118, weq2117, weq2116, weq2115, weq2114, weq2113, weq2112, weq2111, weq2110, weq2109, weq2108, weq2107, weq2106, weq2105, weq2104, weq2103, weq2102, weq2101, weq2100, weq2099, weq2098, weq2097, weq2096, weq2095, weq2094, weq2093, weq2092, weq2091, weq2090, weq2089, weq2088, weq2087, weq2086, weq2085, weq2084, weq2083, weq2082, weq2081, weq2080, weq2079, weq2078, weq2077, weq2076, weq2075, weq2074, weq2073, weq2072, weq2071, weq2070, weq2069, weq2068, weq2067, weq2066, weq2065, weq2064, weq2063, weq2062, weq2061, weq2060, weq2059, weq2058, weq2057, weq2056, weq2055, weq2054, weq2053, weq2052, weq2051, weq2050, weq2049, weq2048, weq2047, weq2046, weq2045, weq2044, weq2043, weq2042, weq2041, weq2040, weq2039, weq2038, weq2037, weq2036, weq2035, weq2034, weq2033, weq2032, weq2031, weq2030, weq2029, weq2028, weq2027, weq2026, weq2025, weq2024, weq2023, weq2022, weq2021, weq2020, weq2019, weq2018, weq2017, weq2016, weq2015, weq2014, weq2013, weq2012, weq2011, weq2010, weq2009, weq2008, weq2007, weq2006, weq2005, weq2004, weq2003, weq2002, weq2001, weq2000, weq1999, weq1998, weq1997, weq1996, weq1995, weq1994, weq1993, weq1992, weq1991, weq1990, weq1989, weq1988, weq1987, weq1986, weq1985, weq1984, weq1983, weq1982, weq1981, weq1980, weq1979, weq1978, weq1977, weq1976, weq1975, weq1974, weq1973, weq1972, weq1971, weq1970, weq1969, weq1968, weq1967, weq1966, weq1965, weq1964, weq1963, weq1962, weq1961, weq1960, weq1959, weq1958, weq1957, weq1956, weq1955, weq1954, weq1953, weq1952, weq1951, weq1950, weq1949, weq1948, weq1947, weq1946, weq1945, weq1944, weq1943, weq1942, weq1941, weq1940, weq1939, weq1938, weq1937, weq1936, weq1935, weq1934, weq1933, weq1932, weq1931, weq1930, weq1929, weq1928, weq1927, weq1926, weq1925, weq1924, weq1923, weq1922, weq1921, weq1920, weq1919, weq1918, weq1917, weq1916, weq1915, weq1914, weq1913, weq1912, weq1911, weq1910, weq1909, weq1908, weq1907, weq1906, weq1905, weq1904, weq1903, weq1902, weq1901, weq1900, weq1899, weq1898, weq1897, weq1896, weq1895, weq1894, weq1893, weq1892, weq1891, weq1890, weq1889, weq1888, weq1887, weq1886, weq1885, weq1884, weq1883, weq1882, weq1881, weq1880, weq1879, weq1878, weq1877, weq1876, weq1875, weq1874, weq1873, weq1872, weq1871, weq1870, weq1869, weq1868, weq1867, weq1866, weq1865, weq1864, weq1863, weq1862, weq1861, weq1860, weq1859, weq1858, weq1857, weq1856, weq1855, weq1854, weq1853, weq1852, weq1851, weq1850, weq1849, weq1848, weq1847, weq1846, weq1845, weq1844, weq1843, weq1842, weq1841, weq1840, weq1839, weq1838, weq1837, weq1836, weq1835, weq1834, weq1833, weq1832, weq1831, weq1830, weq1829, weq1828, weq1827, weq1826, weq1825, weq1824, weq1823, weq1822, weq1821, weq1820, weq1819, weq1818, weq1817, weq1816, weq1815, weq1814, weq1813, weq1812, weq1811, weq1810, weq1809, weq1808, weq1807, weq1806, weq1805, weq1804, weq1803, weq1802, weq1801, weq1800, weq1799, weq1798, weq1797, weq1796, weq1795, weq1794, weq1793, weq1792, weq1791, weq1790, weq1789, weq1788, weq1787, weq1786, weq1785, weq1784, weq1783, weq1782, weq1781, weq1780, weq1779, weq1778, weq1777, weq1776, weq1775, weq1774, weq1773, weq1772, weq1771, weq1770, weq1769, weq1768, weq1767, weq1766, weq1765, weq1764, weq1763, weq1762, weq1761, weq1760, weq1759, weq1758, weq1757, weq1756, weq1755, weq1754, weq1753, weq1752, weq1751, weq1750, weq1749, weq1748, weq1747, weq1746, weq1745, weq1744, weq1743, weq1742, weq1741, weq1740, weq1739, weq1738, weq1737, weq1736, weq1735, weq1734, weq1733, weq1732, weq1731, weq1730, weq1729, weq1728, weq1727, weq1726, weq1725, weq1724, weq1723, weq1722, weq1721, weq1720, weq1719, weq1718, weq1717, weq1716, weq1715, weq1714, weq1713, weq1712, weq1711, weq1710, weq1709, weq1708, weq1707, weq1706, weq1705, weq1704, weq1703, weq1702, weq1701, weq1700, weq1699, weq1698, weq1697, weq1696, weq1695, weq1694, weq1693, weq1692, weq1691, weq1690, weq1689, weq1688, weq1687, weq1686, weq1685, weq1684, weq1683, weq1682, weq1681, weq1680, weq1679, weq1678, weq1677, weq1676, weq1675, weq1674, weq1673, weq1672, weq1671, weq1670, weq1669, weq1668, weq1667, weq1666, weq1665, weq1664, weq1663, weq1662, weq1661, weq1660, weq1659, weq1658, weq1657, weq1656, weq1655, weq1654, weq1653, weq1652, weq1651, weq1650, weq1649, weq1648, weq1647, weq1646, weq1645, weq1644, weq1643, weq1642, weq1641, weq1640, weq1639, weq1638, weq1637, weq1636, weq1635, weq1634, weq1633, weq1632, weq1631, weq1630, weq1629, weq1628, weq1627, weq1626, weq1625, weq1624, weq1623, weq1622, weq1621, weq1620, weq1619, weq1618, weq1617, weq1616, weq1615, weq1614, weq1613, weq1612, weq1611, weq1610, weq1609, weq1608, weq1607, weq1606, weq1605, weq1604, weq1603, weq1602, weq1601, weq1600, weq1599, weq1598, weq1597, weq1596, weq1595, weq1594, weq1593, weq1592, weq1591, weq1590, weq1589, weq1588, weq1587, weq1586, weq1585, weq1584, weq1583, weq1582, weq1581, weq1580, weq1579, weq1578, weq1577, weq1576, weq1575, weq1574, weq1573, weq1572, weq1571, weq1570, weq1569, weq1568, weq1567, weq1566, weq1565, weq1564, weq1563, weq1562, weq1561, weq1560, weq1559, weq1558, weq1557, weq1556, weq1555, weq1554, weq1553, weq1552, weq1551, weq1550, weq1549, weq1548, weq1547, weq1546, weq1545, weq1544, weq1543, weq1542, weq1541, weq1540, weq1539, weq1538, weq1537, weq1536, weq1535, weq1534, weq1533, weq1532, weq1531, weq1530, weq1529, weq1528, weq1527, weq1526, weq1525, weq1524, weq1523, weq1522, weq1521, weq1520, weq1519, weq1518, weq1517, weq1516, weq1515, weq1514, weq1513, weq1512, weq1511, weq1510, weq1509, weq1508, weq1507, weq1506, weq1505, weq1504, weq1503, weq1502, weq1501, weq1500, weq1499, weq1498, weq1497, weq1496, weq1495, weq1494, weq1493, weq1492, weq1491, weq1490, weq1489, weq1488, weq1487, weq1486, weq1485, weq1484, weq1483, weq1482, weq1481, weq1480, weq1479, weq1478, weq1477, weq1476, weq1475, weq1474, weq1473, weq1472, weq1471, weq1470, weq1469, weq1468, weq1467, weq1466, weq1465, weq1464, weq1463, weq1462, weq1461, weq1460, weq1459, weq1458, weq1457, weq1456, weq1455, weq1454, weq1453, weq1452, weq1451, weq1450, weq1449, weq1448, weq1447, weq1446, weq1445, weq1444, weq1443, weq1442, weq1441, weq1440, weq1439, weq1438, weq1437, weq1436, weq1435, weq1434, weq1433, weq1432, weq1431, weq1430, weq1429, weq1428, weq1427, weq1426, weq1425, weq1424, weq1423, weq1422, weq1421, weq1420, weq1419, weq1418, weq1417, weq1416, weq1415, weq1414, weq1413, weq1412, weq1411, weq1410, weq1409, weq1408, weq1407, weq1406, weq1405, weq1404, weq1403, weq1402, weq1401, weq1400, weq1399, weq1398, weq1397, weq1396, weq1395, weq1394, weq1393, weq1392, weq1391, weq1390, weq1389, weq1388, weq1387, weq1386, weq1385, weq1384, weq1383, weq1382, weq1381, weq1380, weq1379, weq1378, weq1377, weq1376, weq1375, weq1374, weq1373, weq1372, weq1371, weq1370, weq1369, weq1368, weq1367, weq1366, weq1365, weq1364, weq1363, weq1362, weq1361, weq1360, weq1359, weq1358, weq1357, weq1356, weq1355, weq1354, weq1353, weq1352, weq1351, weq1350, weq1349, weq1348, weq1347, weq1346, weq1345, weq1344, weq1343, weq1342, weq1341, weq1340, weq1339, weq1338, weq1337, weq1336, weq1335, weq1334, weq1333, weq1332, weq1331, weq1330, weq1329, weq1328, weq1327, weq1326, weq1325, weq1324, weq1323, weq1322, weq1321, weq1320, weq1319, weq1318, weq1317, weq1316, weq1315, weq1314, weq1313, weq1312, weq1311, weq1310, weq1309, weq1308, weq1307, weq1306, weq1305, weq1304, weq1303, weq1302, weq1301, weq1300, weq1299, weq1298, weq1297, weq1296, weq1295, weq1294, weq1293, weq1292, weq1291, weq1290, weq1289, weq1288, weq1287, weq1286, weq1285, weq1284, weq1283, weq1282, weq1281, weq1280, weq1279, weq1278, weq1277, weq1276, weq1275, weq1274, weq1273, weq1272, weq1271, weq1270, weq1269, weq1268, weq1267, weq1266, weq1265, weq1264, weq1263, weq1262, weq1261, weq1260, weq1259, weq1258, weq1257, weq1256, weq1255, weq1254, weq1253, weq1252, weq1251, weq1250, weq1249, weq1248, weq1247, weq1246, weq1245, weq1244, weq1243, weq1242, weq1241, weq1240, weq1239, weq1238, weq1237, weq1236, weq1235, weq1234, weq1233, weq1232, weq1231, weq1230, weq1229, weq1228, weq1227, weq1226, weq1225, weq1224, weq1223, weq1222, weq1221, weq1220, weq1219, weq1218, weq1217, weq1216, weq1215, weq1214, weq1213, weq1212, weq1211, weq1210, weq1209, weq1208, weq1207, weq1206, weq1205, weq1204, weq1203, weq1202, weq1201, weq1200, weq1199, weq1198, weq1197, weq1196, weq1195, weq1194, weq1193, weq1192, weq1191, weq1190, weq1189, weq1188, weq1187, weq1186, weq1185, weq1184, weq1183, weq1182, weq1181, weq1180, weq1179, weq1178, weq1177, weq1176, weq1175, weq1174, weq1173, weq1172, weq1171, weq1170, weq1169, weq1168, weq1167, weq1166, weq1165, weq1164, weq1163, weq1162, weq1161, weq1160, weq1159, weq1158, weq1157, weq1156, weq1155, weq1154, weq1153, weq1152, weq1151, weq1150, weq1149, weq1148, weq1147, weq1146, weq1145, weq1144, weq1143, weq1142, weq1141, weq1140, weq1139, weq1138, weq1137, weq1136, weq1135, weq1134, weq1133, weq1132, weq1131, weq1130, weq1129, weq1128, weq1127, weq1126, weq1125, weq1124, weq1123, weq1122, weq1121, weq1120, weq1119, weq1118, weq1117, weq1116, weq1115, weq1114, weq1113, weq1112, weq1111, weq1110, weq1109, weq1108, weq1107, weq1106, weq1105, weq1104, weq1103, weq1102, weq1101, weq1100, weq1099, weq1098, weq1097, weq1096, weq1095, weq1094, weq1093, weq1092, weq1091, weq1090, weq1089, weq1088, weq1087, weq1086, weq1085, weq1084, weq1083, weq1082, weq1081, weq1080, weq1079, weq1078, weq1077, weq1076, weq1075, weq1074, weq1073, weq1072, weq1071, weq1070, weq1069, weq1068, weq1067, weq1066, weq1065, weq1064, weq1063, weq1062, weq1061, weq1060, weq1059, weq1058, weq1057, weq1056, weq1055, weq1054, weq1053, weq1052, weq1051, weq1050, weq1049, weq1048, weq1047, weq1046, weq1045, weq1044, weq1043, weq1042, weq1041, weq1040, weq1039, weq1038, weq1037, weq1036, weq1035, weq1034, weq1033, weq1032, weq1031, weq1030, weq1029, weq1028, weq1027, weq1026, weq1025, weq1024, weq1023, weq1022, weq1021, weq1020, weq1019, weq1018, weq1017, weq1016, weq1015, weq1014, weq1013, weq1012, weq1011, weq1010, weq1009, weq1008, weq1007, weq1006, weq1005, weq1004, weq1003, weq1002, weq1001, weq1000, weq999, weq998, weq997, weq996, weq995, weq994, weq993, weq992, weq991, weq990, weq989, weq988, weq987, weq986, weq985, weq984, weq983, weq982, weq981, weq980, weq979, weq978, weq977, weq976, weq975, weq974, weq973, weq972, weq971, weq970, weq969, weq968, weq967, weq966, weq965, weq964, weq963, weq962, weq961, weq960, weq959, weq958, weq957, weq956, weq955, weq954, weq953, weq952, weq951, weq950, weq949, weq948, weq947, weq946, weq945, weq944, weq943, weq942, weq941, weq940, weq939, weq938, weq937, weq936, weq935, weq934, weq933, weq932, weq931, weq930, weq929, weq928, weq927, weq926, weq925, weq924, weq923, weq922, weq921, weq920, weq919, weq918, weq917, weq916, weq915, weq914, weq913, weq912, weq911, weq910, weq909, weq908, weq907, weq906, weq905, weq904, weq903, weq902, weq901, weq900, weq899, weq898, weq897, weq896, weq895, weq894, weq893, weq892, weq891, weq890, weq889, weq888, weq887, weq886, weq885, weq884, weq883, weq882, weq881, weq880, weq879, weq878, weq877, weq876, weq875, weq874, weq873, weq872, weq871, weq870, weq869, weq868, weq867, weq866, weq865, weq864, weq863, weq862, weq861, weq860, weq859, weq858, weq857, weq856, weq855, weq854, weq853, weq852, weq851, weq850, weq849, weq848, weq847, weq846, weq845, weq844, weq843, weq842, weq841, weq840, weq839, weq838, weq837, weq836, weq835, weq834, weq833, weq832, weq831, weq830, weq829, weq828, weq827, weq826, weq825, weq824, weq823, weq822, weq821, weq820, weq819, weq818, weq817, weq816, weq815, weq814, weq813, weq812, weq811, weq810, weq809, weq808, weq807, weq806, weq805, weq804, weq803, weq802, weq801, weq800, weq799, weq798, weq797, weq796, weq795, weq794, weq793, weq792, weq791, weq790, weq789, weq788, weq787, weq786, weq785, weq784, weq783, weq782, weq781, weq780, weq779, weq778, weq777, weq776, weq775, weq774, weq773, weq772, weq771, weq770, weq769, weq768, weq767, weq766, weq765, weq764, weq763, weq762, weq761, weq760, weq759, weq758, weq757, weq756, weq755, weq754, weq753, weq752, weq751, weq750, weq749, weq748, weq747, weq746, weq745, weq744, weq743, weq742, weq741, weq740, weq739, weq738, weq737, weq736, weq735, weq734, weq733, weq732, weq731, weq730, weq729, weq728, weq727, weq726, weq725, weq724, weq723, weq722, weq721, weq720, weq719, weq718, weq717, weq716, weq715, weq714, weq713, weq712, weq711, weq710, weq709, weq708, weq707, weq706, weq705, weq704, weq703, weq702, weq701, weq700, weq699, weq698, weq697, weq696, weq695, weq694, weq693, weq692, weq691, weq690, weq689, weq688, weq687, weq686, weq685, weq684, weq683, weq682, weq681, weq680, weq679, weq678, weq677, weq676, weq675, weq674, weq673, weq672, weq671, weq670, weq669, weq668, weq667, weq666, weq665, weq664, weq663, weq662, weq661, weq660, weq659, weq658, weq657, weq656, weq655, weq654, weq653, weq652, weq651, weq650, weq649, weq648, weq647, weq646, weq645, weq644, weq643, weq642, weq641, weq640, weq639, weq638, weq637, weq636, weq635, weq634, weq633, weq632, weq631, weq630, weq629, weq628, weq627, weq626, weq625, weq624, weq623, weq622, weq621, weq620, weq619, weq618, weq617, weq616, weq615, weq614, weq613, weq612, weq611, weq610, weq609, weq608, weq607, weq606, weq605, weq604, weq603, weq602, weq601, weq600, weq599, weq598, weq597, weq596, weq595, weq594, weq593, weq592, weq591, weq590, weq589, weq588, weq587, weq586, weq585, weq584, weq583, weq582, weq581, weq580, weq579, weq578, weq577, weq576, weq575, weq574, weq573, weq572, weq571, weq570, weq569, weq568, weq567, weq566, weq565, weq564, weq563, weq562, weq561, weq560, weq559, weq558, weq557, weq556, weq555, weq554, weq553, weq552, weq551, weq550, weq549, weq548, weq547, weq546, weq545, weq544, weq543, weq542, weq541, weq540, weq539, weq538, weq537, weq536, weq535, weq534, weq533, weq532, weq531, weq530, weq529, weq528, weq527, weq526, weq525, weq524, weq523, weq522, weq521, weq520, weq519, weq518, weq517, weq516, weq515, weq514, weq513, weq512, weq511, weq510, weq509, weq508, weq507, weq506, weq505, weq504, weq503, weq502, weq501, weq500, weq499, weq498, weq497, weq496, weq495, weq494, weq493, weq492, weq491, weq490, weq489, weq488, weq487, weq486, weq485, weq484, weq483, weq482, weq481, weq480, weq479, weq478, weq477, weq476, weq475, weq474, weq473, weq472, weq471, weq470, weq469, weq468, weq467, weq466, weq465, weq464, weq463, weq462, weq461, weq460, weq459, weq458, weq457, weq456, weq455, weq454, weq453, weq452, weq451, weq450, weq449, weq448, weq447, weq446, weq445, weq444, weq443, weq442, weq441, weq440, weq439, weq438, weq437, weq436, weq435, weq434, weq433, weq432, weq431, weq430, weq429, weq428, weq427, weq426, weq425, weq424, weq423, weq422, weq421, weq420, weq419, weq418, weq417, weq416, weq415, weq414, weq413, weq412, weq411, weq410, weq409, weq408, weq407, weq406, weq405, weq404, weq403, weq402, weq401, weq400, weq399, weq398, weq397, weq396, weq395, weq394, weq393, weq392, weq391, weq390, weq389, weq388, weq387, weq386, weq385, weq384, weq383, weq382, weq381, weq380, weq379, weq378, weq377, weq376, weq375, weq374, weq373, weq372, weq371, weq370, weq369, weq368, weq367, weq366, weq365, weq364, weq363, weq362, weq361, weq360, weq359, weq358, weq357, weq356, weq355, weq354, weq353, weq352, weq351, weq350, weq349, weq348, weq347, weq346, weq345, weq344, weq343, weq342, weq341, weq340, weq339, weq338, weq337, weq336, weq335, weq334, weq333, weq332, weq331, weq330, weq329, weq328, weq327, weq326, weq325, weq324, weq323, weq322, weq321, weq320, weq319, weq318, weq317, weq316, weq315, weq314, weq313, weq312, weq311, weq310, weq309, weq308, weq307, weq306, weq305, weq304, weq303, weq302, weq301, weq300, weq299, weq298, weq297, weq296, weq295, weq294, weq293, weq292, weq291, weq290, weq289, weq288, weq287, weq286, weq285, weq284, weq283, weq282, weq281, weq280, weq279, weq278, weq277, weq276, weq275, weq274, weq273, weq272, weq271, weq270, weq269, weq268, weq267, weq266, weq265, weq264, weq263, weq262, weq261, weq260, weq259, weq258, weq257, weq256, weq255, weq254, weq253, weq252, weq251, weq250, weq249, weq248, weq247, weq246, weq245, weq244, weq243, weq242, weq241, weq240, weq239, weq238, weq237, weq236, weq235, weq234, weq233, weq232, weq231, weq230, weq229, weq228, weq227, weq226, weq225, weq224, weq223, weq222, weq221, weq220, weq219, weq218, weq217, weq216, weq215, weq214, weq213, weq212, weq211, weq210, weq209, weq208, weq207, weq206, weq205, weq204, weq203, weq202, weq201, weq200, weq199, weq198, weq197, weq196, weq195, weq194, weq193, weq192, weq191, weq190, weq189, weq188, weq187, weq186, weq185, weq184, weq183, weq182, weq181, weq180, weq179, weq178, weq177, weq176, weq175, weq174, weq173, weq172, weq171, weq170, weq169, weq168, weq167, weq166, weq165, weq164, weq163, weq162, weq161, weq160, weq159, weq158, weq157, weq156, weq155, weq154, weq153, weq152, weq151, weq150, weq149, weq148, weq147, weq146, weq145, weq144, weq143, weq142, weq141, weq140, weq139, weq138, weq137, weq136, weq135, weq134, weq133, weq132, weq131, weq130, weq129, weq128, weq127, weq126, weq125, weq124, weq123, weq122, weq121, weq120, weq119, weq118, weq117, weq116, weq115, weq114, weq113, weq112, weq111, weq110, weq109, weq108, weq107, weq106, weq105, weq104, weq103, weq102, weq101, weq100, weq99, weq98, weq97, weq96, weq95, weq94, weq93, weq92, weq91, weq90, weq89, weq88, weq87, weq86, weq85, weq84, weq83, weq82, weq81, weq80, weq79, weq78, weq77, weq76, weq75, weq74, weq73, weq72, weq71, weq70, weq69, weq68, weq67, weq66, weq65, weq64, weq63, weq62, weq61, weq60, weq59, weq58, weq57, weq56, weq55, weq54, weq53, weq52, weq51, weq50, weq49, weq48, weq47, weq46, weq45, weq44, weq43, weq42, weq41, weq40, weq39, weq38, weq37, weq36, weq35, weq34, weq33, weq32, weq31, weq30, weq29, weq28, weq27, weq26, weq25, weq24, weq23, weq22, weq21, weq20, weq19, weq18, weq17, weq16, weq15, weq14, weq13, weq12, weq11, weq10, weq9, weq8, weq7, weq6, weq5, weq4, weq3, weq2, weq1, weq0};


endmodule