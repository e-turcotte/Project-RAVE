module decode_TOP;
    //instantiate queued latches here? or take in as input?

    

endmodule