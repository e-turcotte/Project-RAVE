module brlogic_t();

endmodule