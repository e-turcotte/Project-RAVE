module prefix_lut(
    input [7:0] prefix1,
    input [7:0] prefix2,
    input [7:0] prefix3,
    output [1:0] num_prefixes,
    output is_rep,
    output is_seg_override,
    output is_opsiz_override
    );

    //compare each prefix to the known prefixes in lookup table
    
    


endmodule