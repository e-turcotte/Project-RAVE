module outputAlign(
    
);

endmodule