module execute_TOP(

);


endmodule 