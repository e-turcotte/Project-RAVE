module instruction_length(
    input wire [11:0] in,
    output wire [7:0] out
);
    wire [11:0] buffered_input;
    wire [7:0] wire0, wire1, wire2, wire3, wire4, wire5, wire6, wire7, wire8, wire9, wire10, wire11, wire12, wire13, wire14, wire15, wire16, wire17, wire18, wire19, wire20, wire21, wire22, wire23, wire24, wire25, wire26, wire27, wire28, wire29, wire30, wire31, wire32, wire33, wire34, wire35, wire36, wire37, wire38, wire39, wire40, wire41, wire42, wire43, wire44, wire45, wire46, wire47, wire48, wire49, wire50, wire51, wire52, wire53, wire54, wire55, wire56, wire57, wire58, wire59, wire60, wire61, wire62, wire63, wire64, wire65, wire66, wire67, wire68, wire69, wire70, wire71, wire72, wire73, wire74, wire75, wire76, wire77, wire78, wire79, wire80, wire81, wire82, wire83, wire84, wire85, wire86, wire87, wire88, wire89, wire90, wire91, wire92, wire93, wire94, wire95, wire96, wire97, wire98, wire99, wire100, wire101, wire102, wire103, wire104, wire105, wire106, wire107, wire108, wire109, wire110, wire111, wire112, wire113, wire114, wire115, wire116, wire117, wire118, wire119, wire120, wire121, wire122, wire123, wire124, wire125, wire126, wire127, wire128, wire129, wire130, wire131, wire132, wire133, wire134, wire135, wire136, wire137, wire138, wire139, wire140, wire141, wire142, wire143, wire144, wire145, wire146, wire147, wire148, wire149, wire150, wire151, wire152, wire153, wire154, wire155, wire156, wire157, wire158, wire159, wire160, wire161, wire162, wire163, wire164, wire165, wire166, wire167, wire168, wire169, wire170, wire171, wire172, wire173, wire174, wire175, wire176, wire177, wire178, wire179, wire180, wire181, wire182, wire183, wire184, wire185, wire186, wire187, wire188, wire189, wire190, wire191, wire192, wire193, wire194, wire195, wire196, wire197, wire198, wire199, wire200, wire201, wire202, wire203, wire204, wire205, wire206, wire207, wire208, wire209, wire210, wire211, wire212, wire213, wire214, wire215, wire216, wire217, wire218, wire219, wire220, wire221, wire222, wire223, wire224, wire225, wire226, wire227, wire228, wire229, wire230, wire231, wire232, wire233, wire234, wire235, wire236, wire237, wire238, wire239, wire240, wire241, wire242, wire243, wire244, wire245, wire246, wire247, wire248, wire249, wire250, wire251, wire252, wire253, wire254, wire255, wire256, wire257, wire258, wire259, wire260, wire261, wire262, wire263, wire264, wire265, wire266, wire267, wire268, wire269, wire270, wire271, wire272, wire273, wire274, wire275, wire276, wire277, wire278, wire279, wire280, wire281, wire282, wire283, wire284, wire285, wire286, wire287, wire288, wire289, wire290, wire291, wire292, wire293, wire294, wire295, wire296, wire297, wire298, wire299, wire300, wire301, wire302, wire303, wire304, wire305, wire306, wire307, wire308, wire309, wire310, wire311, wire312, wire313, wire314, wire315, wire316, wire317, wire318, wire319, wire320, wire321, wire322, wire323, wire324, wire325, wire326, wire327, wire328, wire329, wire330, wire331, wire332, wire333, wire334, wire335, wire336, wire337, wire338, wire339, wire340, wire341, wire342, wire343, wire344, wire345, wire346, wire347, wire348, wire349, wire350, wire351, wire352, wire353, wire354, wire355, wire356, wire357, wire358, wire359, wire360, wire361, wire362, wire363, wire364, wire365, wire366, wire367, wire368, wire369, wire370, wire371, wire372, wire373, wire374, wire375, wire376, wire377, wire378, wire379, wire380, wire381, wire382, wire383, wire384, wire385, wire386, wire387, wire388, wire389, wire390, wire391, wire392, wire393, wire394, wire395, wire396, wire397, wire398, wire399, wire400, wire401, wire402, wire403, wire404, wire405, wire406, wire407, wire408, wire409, wire410, wire411, wire412, wire413, wire414, wire415, wire416, wire417, wire418, wire419, wire420, wire421, wire422, wire423, wire424, wire425, wire426, wire427, wire428, wire429, wire430, wire431, wire432, wire433, wire434, wire435, wire436, wire437, wire438, wire439, wire440, wire441, wire442, wire443, wire444, wire445, wire446, wire447, wire448, wire449, wire450, wire451, wire452, wire453, wire454, wire455, wire456, wire457, wire458, wire459, wire460, wire461, wire462, wire463, wire464, wire465, wire466, wire467, wire468, wire469, wire470, wire471, wire472, wire473, wire474, wire475, wire476, wire477, wire478, wire479, wire480, wire481, wire482, wire483, wire484, wire485, wire486, wire487, wire488, wire489, wire490, wire491, wire492, wire493, wire494, wire495, wire496, wire497, wire498, wire499, wire500, wire501, wire502, wire503, wire504, wire505, wire506, wire507, wire508, wire509, wire510, wire511, wire512, wire513, wire514, wire515, wire516, wire517, wire518, wire519, wire520, wire521, wire522, wire523, wire524, wire525, wire526, wire527, wire528, wire529, wire530, wire531, wire532, wire533, wire534, wire535, wire536, wire537, wire538, wire539, wire540, wire541, wire542, wire543, wire544, wire545, wire546, wire547, wire548, wire549, wire550, wire551, wire552, wire553, wire554, wire555, wire556, wire557, wire558, wire559, wire560, wire561, wire562, wire563, wire564, wire565, wire566, wire567, wire568, wire569, wire570, wire571, wire572, wire573, wire574, wire575, wire576, wire577, wire578, wire579, wire580, wire581, wire582, wire583, wire584, wire585, wire586, wire587, wire588, wire589, wire590, wire591, wire592, wire593, wire594, wire595, wire596, wire597, wire598, wire599, wire600, wire601, wire602, wire603, wire604, wire605, wire606, wire607, wire608, wire609, wire610, wire611, wire612, wire613, wire614, wire615, wire616, wire617, wire618, wire619, wire620, wire621, wire622, wire623, wire624, wire625, wire626, wire627, wire628, wire629, wire630, wire631, wire632, wire633, wire634, wire635, wire636, wire637, wire638, wire639, wire640, wire641, wire642, wire643, wire644, wire645, wire646, wire647, wire648, wire649, wire650, wire651, wire652, wire653, wire654, wire655, wire656, wire657, wire658, wire659, wire660, wire661, wire662, wire663, wire664, wire665, wire666, wire667, wire668, wire669, wire670, wire671, wire672, wire673, wire674, wire675, wire676, wire677, wire678, wire679, wire680, wire681, wire682, wire683, wire684, wire685, wire686, wire687, wire688, wire689, wire690, wire691, wire692, wire693, wire694, wire695, wire696, wire697, wire698, wire699, wire700, wire701, wire702, wire703, wire704, wire705, wire706, wire707, wire708, wire709, wire710, wire711, wire712, wire713, wire714, wire715, wire716, wire717, wire718, wire719, wire720, wire721, wire722, wire723, wire724, wire725, wire726, wire727, wire728, wire729, wire730, wire731, wire732, wire733, wire734, wire735, wire736, wire737, wire738, wire739, wire740, wire741, wire742, wire743, wire744, wire745, wire746, wire747, wire748, wire749, wire750, wire751, wire752, wire753, wire754, wire755, wire756, wire757, wire758, wire759, wire760, wire761, wire762, wire763, wire764, wire765, wire766, wire767, wire768, wire769, wire770, wire771, wire772, wire773, wire774, wire775, wire776, wire777, wire778, wire779, wire780, wire781, wire782, wire783, wire784, wire785, wire786, wire787, wire788, wire789, wire790, wire791, wire792, wire793, wire794, wire795, wire796, wire797, wire798, wire799, wire800, wire801, wire802, wire803, wire804, wire805, wire806, wire807, wire808, wire809, wire810, wire811, wire812, wire813, wire814, wire815, wire816, wire817, wire818, wire819, wire820, wire821, wire822, wire823, wire824, wire825, wire826, wire827, wire828, wire829, wire830, wire831, wire832, wire833, wire834, wire835, wire836, wire837, wire838, wire839, wire840, wire841, wire842, wire843, wire844, wire845, wire846, wire847, wire848, wire849, wire850, wire851, wire852, wire853, wire854, wire855, wire856, wire857, wire858, wire859, wire860, wire861, wire862, wire863, wire864, wire865, wire866, wire867, wire868, wire869, wire870, wire871, wire872, wire873, wire874, wire875, wire876, wire877, wire878, wire879, wire880, wire881, wire882, wire883, wire884, wire885, wire886, wire887, wire888, wire889, wire890, wire891, wire892, wire893, wire894, wire895, wire896, wire897, wire898, wire899, wire900, wire901, wire902, wire903, wire904, wire905, wire906, wire907, wire908, wire909, wire910, wire911, wire912, wire913, wire914, wire915, wire916, wire917, wire918, wire919, wire920, wire921, wire922, wire923, wire924, wire925, wire926, wire927, wire928, wire929, wire930, wire931, wire932, wire933, wire934, wire935, wire936, wire937, wire938, wire939, wire940, wire941, wire942, wire943, wire944, wire945, wire946, wire947, wire948, wire949, wire950, wire951, wire952, wire953, wire954, wire955, wire956, wire957, wire958, wire959, wire960, wire961, wire962, wire963, wire964, wire965, wire966, wire967, wire968, wire969, wire970, wire971, wire972, wire973, wire974, wire975, wire976, wire977, wire978, wire979, wire980, wire981, wire982, wire983, wire984, wire985, wire986, wire987, wire988, wire989, wire990, wire991, wire992, wire993, wire994, wire995, wire996, wire997, wire998, wire999, wire1000, wire1001, wire1002, wire1003, wire1004, wire1005, wire1006, wire1007, wire1008, wire1009, wire1010, wire1011, wire1012, wire1013, wire1014, wire1015, wire1016, wire1017, wire1018, wire1019, wire1020, wire1021, wire1022, wire1023, wire1024, wire1025, wire1026, wire1027, wire1028, wire1029, wire1030, wire1031, wire1032, wire1033, wire1034, wire1035, wire1036, wire1037, wire1038, wire1039, wire1040, wire1041, wire1042, wire1043, wire1044, wire1045, wire1046, wire1047, wire1048, wire1049, wire1050, wire1051, wire1052, wire1053, wire1054, wire1055, wire1056, wire1057, wire1058, wire1059, wire1060, wire1061, wire1062, wire1063, wire1064, wire1065, wire1066, wire1067, wire1068, wire1069, wire1070, wire1071, wire1072, wire1073, wire1074, wire1075, wire1076, wire1077, wire1078, wire1079, wire1080, wire1081, wire1082, wire1083, wire1084, wire1085, wire1086, wire1087, wire1088, wire1089, wire1090, wire1091, wire1092, wire1093, wire1094, wire1095, wire1096, wire1097, wire1098, wire1099, wire1100, wire1101, wire1102, wire1103, wire1104, wire1105, wire1106, wire1107, wire1108, wire1109, wire1110, wire1111, wire1112, wire1113, wire1114, wire1115, wire1116, wire1117, wire1118, wire1119, wire1120, wire1121, wire1122, wire1123, wire1124, wire1125, wire1126, wire1127, wire1128, wire1129, wire1130, wire1131, wire1132, wire1133, wire1134, wire1135, wire1136, wire1137, wire1138, wire1139, wire1140, wire1141, wire1142, wire1143, wire1144, wire1145, wire1146, wire1147, wire1148, wire1149, wire1150, wire1151, wire1152, wire1153, wire1154, wire1155, wire1156, wire1157, wire1158, wire1159, wire1160, wire1161, wire1162, wire1163, wire1164, wire1165, wire1166, wire1167, wire1168, wire1169, wire1170, wire1171, wire1172, wire1173, wire1174, wire1175, wire1176, wire1177, wire1178, wire1179, wire1180, wire1181, wire1182, wire1183, wire1184, wire1185, wire1186, wire1187, wire1188, wire1189, wire1190, wire1191, wire1192, wire1193, wire1194, wire1195, wire1196, wire1197, wire1198, wire1199, wire1200, wire1201, wire1202, wire1203, wire1204, wire1205, wire1206, wire1207, wire1208, wire1209, wire1210, wire1211, wire1212, wire1213, wire1214, wire1215, wire1216, wire1217, wire1218, wire1219, wire1220, wire1221, wire1222, wire1223, wire1224, wire1225, wire1226, wire1227, wire1228, wire1229, wire1230, wire1231, wire1232, wire1233, wire1234, wire1235, wire1236, wire1237, wire1238, wire1239, wire1240, wire1241, wire1242, wire1243, wire1244, wire1245, wire1246, wire1247, wire1248, wire1249, wire1250, wire1251, wire1252, wire1253, wire1254, wire1255, wire1256, wire1257, wire1258, wire1259, wire1260, wire1261, wire1262, wire1263, wire1264, wire1265, wire1266, wire1267, wire1268, wire1269, wire1270, wire1271, wire1272, wire1273, wire1274, wire1275, wire1276, wire1277, wire1278, wire1279, wire1280, wire1281, wire1282, wire1283, wire1284, wire1285, wire1286, wire1287, wire1288, wire1289, wire1290, wire1291, wire1292, wire1293, wire1294, wire1295, wire1296, wire1297, wire1298, wire1299, wire1300, wire1301, wire1302, wire1303, wire1304, wire1305, wire1306, wire1307, wire1308, wire1309, wire1310, wire1311, wire1312, wire1313, wire1314, wire1315, wire1316, wire1317, wire1318, wire1319, wire1320, wire1321, wire1322, wire1323, wire1324, wire1325, wire1326, wire1327, wire1328, wire1329, wire1330, wire1331, wire1332, wire1333, wire1334, wire1335, wire1336, wire1337, wire1338, wire1339, wire1340, wire1341, wire1342, wire1343, wire1344, wire1345, wire1346, wire1347, wire1348, wire1349, wire1350, wire1351, wire1352, wire1353, wire1354, wire1355, wire1356, wire1357, wire1358, wire1359, wire1360, wire1361, wire1362, wire1363, wire1364, wire1365, wire1366, wire1367, wire1368, wire1369, wire1370, wire1371, wire1372, wire1373, wire1374, wire1375, wire1376, wire1377, wire1378, wire1379, wire1380, wire1381, wire1382, wire1383, wire1384, wire1385, wire1386, wire1387, wire1388, wire1389, wire1390, wire1391, wire1392, wire1393, wire1394, wire1395, wire1396, wire1397, wire1398, wire1399, wire1400, wire1401, wire1402, wire1403, wire1404, wire1405, wire1406, wire1407, wire1408, wire1409, wire1410, wire1411, wire1412, wire1413, wire1414, wire1415, wire1416, wire1417, wire1418, wire1419, wire1420, wire1421, wire1422, wire1423, wire1424, wire1425, wire1426, wire1427, wire1428, wire1429, wire1430, wire1431, wire1432, wire1433, wire1434, wire1435, wire1436, wire1437, wire1438, wire1439, wire1440, wire1441, wire1442, wire1443, wire1444, wire1445, wire1446, wire1447, wire1448, wire1449, wire1450, wire1451, wire1452, wire1453, wire1454, wire1455, wire1456, wire1457, wire1458, wire1459, wire1460, wire1461, wire1462, wire1463, wire1464, wire1465, wire1466, wire1467, wire1468, wire1469, wire1470, wire1471, wire1472, wire1473, wire1474, wire1475, wire1476, wire1477, wire1478, wire1479, wire1480, wire1481, wire1482, wire1483, wire1484, wire1485, wire1486, wire1487, wire1488, wire1489, wire1490, wire1491, wire1492, wire1493, wire1494, wire1495, wire1496, wire1497, wire1498, wire1499, wire1500, wire1501, wire1502, wire1503, wire1504, wire1505, wire1506, wire1507, wire1508, wire1509, wire1510, wire1511, wire1512, wire1513, wire1514, wire1515, wire1516, wire1517, wire1518, wire1519, wire1520, wire1521, wire1522, wire1523, wire1524, wire1525, wire1526, wire1527, wire1528, wire1529, wire1530, wire1531, wire1532, wire1533, wire1534, wire1535, wire1536, wire1537, wire1538, wire1539, wire1540, wire1541, wire1542, wire1543, wire1544, wire1545, wire1546, wire1547, wire1548, wire1549, wire1550, wire1551, wire1552, wire1553, wire1554, wire1555, wire1556, wire1557, wire1558, wire1559, wire1560, wire1561, wire1562, wire1563, wire1564, wire1565, wire1566, wire1567, wire1568, wire1569, wire1570, wire1571, wire1572, wire1573, wire1574, wire1575, wire1576, wire1577, wire1578, wire1579, wire1580, wire1581, wire1582, wire1583, wire1584, wire1585, wire1586, wire1587, wire1588, wire1589, wire1590, wire1591, wire1592, wire1593, wire1594, wire1595, wire1596, wire1597, wire1598, wire1599, wire1600, wire1601, wire1602, wire1603, wire1604, wire1605, wire1606, wire1607, wire1608, wire1609, wire1610, wire1611, wire1612, wire1613, wire1614, wire1615, wire1616, wire1617, wire1618, wire1619, wire1620, wire1621, wire1622, wire1623, wire1624, wire1625, wire1626, wire1627, wire1628, wire1629, wire1630, wire1631, wire1632, wire1633, wire1634, wire1635, wire1636, wire1637, wire1638, wire1639, wire1640, wire1641, wire1642, wire1643, wire1644, wire1645, wire1646, wire1647, wire1648, wire1649, wire1650, wire1651, wire1652, wire1653, wire1654, wire1655, wire1656, wire1657, wire1658, wire1659, wire1660, wire1661, wire1662, wire1663, wire1664, wire1665, wire1666, wire1667, wire1668, wire1669, wire1670, wire1671, wire1672, wire1673, wire1674, wire1675, wire1676, wire1677, wire1678, wire1679, wire1680, wire1681, wire1682, wire1683, wire1684, wire1685, wire1686, wire1687, wire1688, wire1689, wire1690, wire1691, wire1692, wire1693, wire1694, wire1695, wire1696, wire1697, wire1698, wire1699, wire1700, wire1701, wire1702, wire1703, wire1704, wire1705, wire1706, wire1707, wire1708, wire1709, wire1710, wire1711, wire1712, wire1713, wire1714, wire1715, wire1716, wire1717, wire1718, wire1719, wire1720, wire1721, wire1722, wire1723, wire1724, wire1725, wire1726, wire1727, wire1728, wire1729, wire1730, wire1731, wire1732, wire1733, wire1734, wire1735, wire1736, wire1737, wire1738, wire1739, wire1740, wire1741, wire1742, wire1743, wire1744, wire1745, wire1746, wire1747, wire1748, wire1749, wire1750, wire1751, wire1752, wire1753, wire1754, wire1755, wire1756, wire1757, wire1758, wire1759, wire1760, wire1761, wire1762, wire1763, wire1764, wire1765, wire1766, wire1767, wire1768, wire1769, wire1770, wire1771, wire1772, wire1773, wire1774, wire1775, wire1776, wire1777, wire1778, wire1779, wire1780, wire1781, wire1782, wire1783, wire1784, wire1785, wire1786, wire1787, wire1788, wire1789, wire1790, wire1791, wire1792, wire1793, wire1794, wire1795, wire1796, wire1797, wire1798, wire1799, wire1800, wire1801, wire1802, wire1803, wire1804, wire1805, wire1806, wire1807, wire1808, wire1809, wire1810, wire1811, wire1812, wire1813, wire1814, wire1815, wire1816, wire1817, wire1818, wire1819, wire1820, wire1821, wire1822, wire1823, wire1824, wire1825, wire1826, wire1827, wire1828, wire1829, wire1830, wire1831, wire1832, wire1833, wire1834, wire1835, wire1836, wire1837, wire1838, wire1839, wire1840, wire1841, wire1842, wire1843, wire1844, wire1845, wire1846, wire1847, wire1848, wire1849, wire1850, wire1851, wire1852, wire1853, wire1854, wire1855, wire1856, wire1857, wire1858, wire1859, wire1860, wire1861, wire1862, wire1863, wire1864, wire1865, wire1866, wire1867, wire1868, wire1869, wire1870, wire1871, wire1872, wire1873, wire1874, wire1875, wire1876, wire1877, wire1878, wire1879, wire1880, wire1881, wire1882, wire1883, wire1884, wire1885, wire1886, wire1887, wire1888, wire1889, wire1890, wire1891, wire1892, wire1893, wire1894, wire1895, wire1896, wire1897, wire1898, wire1899, wire1900, wire1901, wire1902, wire1903, wire1904, wire1905, wire1906, wire1907, wire1908, wire1909, wire1910, wire1911, wire1912, wire1913, wire1914, wire1915, wire1916, wire1917, wire1918, wire1919, wire1920, wire1921, wire1922, wire1923, wire1924, wire1925, wire1926, wire1927, wire1928, wire1929, wire1930, wire1931, wire1932, wire1933, wire1934, wire1935, wire1936, wire1937, wire1938, wire1939, wire1940, wire1941, wire1942, wire1943, wire1944, wire1945, wire1946, wire1947, wire1948, wire1949, wire1950, wire1951, wire1952, wire1953, wire1954, wire1955, wire1956, wire1957, wire1958, wire1959, wire1960, wire1961, wire1962, wire1963, wire1964, wire1965, wire1966, wire1967, wire1968, wire1969, wire1970, wire1971, wire1972, wire1973, wire1974, wire1975, wire1976, wire1977, wire1978, wire1979, wire1980, wire1981, wire1982, wire1983, wire1984, wire1985, wire1986, wire1987, wire1988, wire1989, wire1990, wire1991, wire1992, wire1993, wire1994, wire1995, wire1996, wire1997, wire1998, wire1999, wire2000, wire2001, wire2002, wire2003, wire2004, wire2005, wire2006, wire2007, wire2008, wire2009, wire2010, wire2011, wire2012, wire2013, wire2014, wire2015, wire2016, wire2017, wire2018, wire2019, wire2020, wire2021, wire2022, wire2023, wire2024, wire2025, wire2026, wire2027, wire2028, wire2029, wire2030, wire2031, wire2032, wire2033, wire2034, wire2035, wire2036, wire2037, wire2038, wire2039, wire2040, wire2041, wire2042, wire2043, wire2044, wire2045, wire2046, wire2047, wire2048, wire2049, wire2050, wire2051, wire2052, wire2053, wire2054, wire2055, wire2056, wire2057, wire2058, wire2059, wire2060, wire2061, wire2062, wire2063, wire2064, wire2065, wire2066, wire2067, wire2068, wire2069, wire2070, wire2071, wire2072, wire2073, wire2074, wire2075, wire2076, wire2077, wire2078, wire2079, wire2080, wire2081, wire2082, wire2083, wire2084, wire2085, wire2086, wire2087, wire2088, wire2089, wire2090, wire2091, wire2092, wire2093, wire2094, wire2095, wire2096, wire2097, wire2098, wire2099, wire2100, wire2101, wire2102, wire2103, wire2104, wire2105, wire2106, wire2107, wire2108, wire2109, wire2110, wire2111, wire2112, wire2113, wire2114, wire2115, wire2116, wire2117, wire2118, wire2119, wire2120, wire2121, wire2122, wire2123, wire2124, wire2125, wire2126, wire2127, wire2128, wire2129, wire2130, wire2131, wire2132, wire2133, wire2134, wire2135, wire2136, wire2137, wire2138, wire2139, wire2140, wire2141, wire2142, wire2143, wire2144, wire2145, wire2146, wire2147, wire2148, wire2149, wire2150, wire2151, wire2152, wire2153, wire2154, wire2155, wire2156, wire2157, wire2158, wire2159, wire2160, wire2161, wire2162, wire2163, wire2164, wire2165, wire2166, wire2167, wire2168, wire2169, wire2170, wire2171, wire2172, wire2173, wire2174, wire2175, wire2176, wire2177, wire2178, wire2179, wire2180, wire2181, wire2182, wire2183, wire2184, wire2185, wire2186, wire2187, wire2188, wire2189, wire2190, wire2191, wire2192, wire2193, wire2194, wire2195, wire2196, wire2197, wire2198, wire2199, wire2200, wire2201, wire2202, wire2203, wire2204, wire2205, wire2206, wire2207, wire2208, wire2209, wire2210, wire2211, wire2212, wire2213, wire2214, wire2215, wire2216, wire2217, wire2218, wire2219, wire2220, wire2221, wire2222, wire2223, wire2224, wire2225, wire2226, wire2227, wire2228, wire2229, wire2230, wire2231, wire2232, wire2233, wire2234, wire2235, wire2236, wire2237, wire2238, wire2239, wire2240, wire2241, wire2242, wire2243, wire2244, wire2245, wire2246, wire2247, wire2248, wire2249, wire2250, wire2251, wire2252, wire2253, wire2254, wire2255, wire2256, wire2257, wire2258, wire2259, wire2260, wire2261, wire2262, wire2263, wire2264, wire2265, wire2266, wire2267, wire2268, wire2269, wire2270, wire2271, wire2272, wire2273, wire2274, wire2275, wire2276, wire2277, wire2278, wire2279, wire2280, wire2281, wire2282, wire2283, wire2284, wire2285, wire2286, wire2287, wire2288, wire2289, wire2290, wire2291, wire2292, wire2293, wire2294, wire2295, wire2296, wire2297, wire2298, wire2299, wire2300, wire2301, wire2302, wire2303, wire2304, wire2305, wire2306, wire2307, wire2308, wire2309, wire2310, wire2311, wire2312, wire2313, wire2314, wire2315, wire2316, wire2317, wire2318, wire2319, wire2320, wire2321, wire2322, wire2323, wire2324, wire2325, wire2326, wire2327, wire2328, wire2329, wire2330, wire2331, wire2332, wire2333, wire2334, wire2335, wire2336, wire2337, wire2338, wire2339, wire2340, wire2341, wire2342, wire2343, wire2344, wire2345, wire2346, wire2347, wire2348, wire2349, wire2350, wire2351, wire2352, wire2353, wire2354, wire2355, wire2356, wire2357, wire2358, wire2359, wire2360, wire2361, wire2362, wire2363, wire2364, wire2365, wire2366, wire2367, wire2368, wire2369, wire2370, wire2371, wire2372, wire2373, wire2374, wire2375, wire2376, wire2377, wire2378, wire2379, wire2380, wire2381, wire2382, wire2383, wire2384, wire2385, wire2386, wire2387, wire2388, wire2389, wire2390, wire2391, wire2392, wire2393, wire2394, wire2395, wire2396, wire2397, wire2398, wire2399, wire2400, wire2401, wire2402, wire2403, wire2404, wire2405, wire2406, wire2407, wire2408, wire2409, wire2410, wire2411, wire2412, wire2413, wire2414, wire2415, wire2416, wire2417, wire2418, wire2419, wire2420, wire2421, wire2422, wire2423, wire2424, wire2425, wire2426, wire2427, wire2428, wire2429, wire2430, wire2431, wire2432, wire2433, wire2434, wire2435, wire2436, wire2437, wire2438, wire2439, wire2440, wire2441, wire2442, wire2443, wire2444, wire2445, wire2446, wire2447, wire2448, wire2449, wire2450, wire2451, wire2452, wire2453, wire2454, wire2455, wire2456, wire2457, wire2458, wire2459, wire2460, wire2461, wire2462, wire2463, wire2464, wire2465, wire2466, wire2467, wire2468, wire2469, wire2470, wire2471, wire2472, wire2473, wire2474, wire2475, wire2476, wire2477, wire2478, wire2479, wire2480, wire2481, wire2482, wire2483, wire2484, wire2485, wire2486, wire2487, wire2488, wire2489, wire2490, wire2491, wire2492, wire2493, wire2494, wire2495, wire2496, wire2497, wire2498, wire2499, wire2500, wire2501, wire2502, wire2503, wire2504, wire2505, wire2506, wire2507, wire2508, wire2509, wire2510, wire2511, wire2512, wire2513, wire2514, wire2515, wire2516, wire2517, wire2518, wire2519, wire2520, wire2521, wire2522, wire2523, wire2524, wire2525, wire2526, wire2527, wire2528, wire2529, wire2530, wire2531, wire2532, wire2533, wire2534, wire2535, wire2536, wire2537, wire2538, wire2539, wire2540, wire2541, wire2542, wire2543, wire2544, wire2545, wire2546, wire2547, wire2548, wire2549, wire2550, wire2551, wire2552, wire2553, wire2554, wire2555, wire2556, wire2557, wire2558, wire2559, wire2560, wire2561, wire2562, wire2563, wire2564, wire2565, wire2566, wire2567, wire2568, wire2569, wire2570, wire2571, wire2572, wire2573, wire2574, wire2575, wire2576, wire2577, wire2578, wire2579, wire2580, wire2581, wire2582, wire2583, wire2584, wire2585, wire2586, wire2587, wire2588, wire2589, wire2590, wire2591, wire2592, wire2593, wire2594, wire2595, wire2596, wire2597, wire2598, wire2599, wire2600, wire2601, wire2602, wire2603, wire2604, wire2605, wire2606, wire2607, wire2608, wire2609, wire2610, wire2611, wire2612, wire2613, wire2614, wire2615, wire2616, wire2617, wire2618, wire2619, wire2620, wire2621, wire2622, wire2623, wire2624, wire2625, wire2626, wire2627, wire2628, wire2629, wire2630, wire2631, wire2632, wire2633, wire2634, wire2635, wire2636, wire2637, wire2638, wire2639, wire2640, wire2641, wire2642, wire2643, wire2644, wire2645, wire2646, wire2647, wire2648, wire2649, wire2650, wire2651, wire2652, wire2653, wire2654, wire2655, wire2656, wire2657, wire2658, wire2659, wire2660, wire2661, wire2662, wire2663, wire2664, wire2665, wire2666, wire2667, wire2668, wire2669, wire2670, wire2671, wire2672, wire2673, wire2674, wire2675, wire2676, wire2677, wire2678, wire2679, wire2680, wire2681, wire2682, wire2683, wire2684, wire2685, wire2686, wire2687, wire2688, wire2689, wire2690, wire2691, wire2692, wire2693, wire2694, wire2695, wire2696, wire2697, wire2698, wire2699, wire2700, wire2701, wire2702, wire2703, wire2704, wire2705, wire2706, wire2707, wire2708, wire2709, wire2710, wire2711, wire2712, wire2713, wire2714, wire2715, wire2716, wire2717, wire2718, wire2719, wire2720, wire2721, wire2722, wire2723, wire2724, wire2725, wire2726, wire2727, wire2728, wire2729, wire2730, wire2731, wire2732, wire2733, wire2734, wire2735, wire2736, wire2737, wire2738, wire2739, wire2740, wire2741, wire2742, wire2743, wire2744, wire2745, wire2746, wire2747, wire2748, wire2749, wire2750, wire2751, wire2752, wire2753, wire2754, wire2755, wire2756, wire2757, wire2758, wire2759, wire2760, wire2761, wire2762, wire2763, wire2764, wire2765, wire2766, wire2767, wire2768, wire2769, wire2770, wire2771, wire2772, wire2773, wire2774, wire2775, wire2776, wire2777, wire2778, wire2779, wire2780, wire2781, wire2782, wire2783, wire2784, wire2785, wire2786, wire2787, wire2788, wire2789, wire2790, wire2791, wire2792, wire2793, wire2794, wire2795, wire2796, wire2797, wire2798, wire2799, wire2800, wire2801, wire2802, wire2803, wire2804, wire2805, wire2806, wire2807, wire2808, wire2809, wire2810, wire2811, wire2812, wire2813, wire2814, wire2815, wire2816, wire2817, wire2818, wire2819, wire2820, wire2821, wire2822, wire2823, wire2824, wire2825, wire2826, wire2827, wire2828, wire2829, wire2830, wire2831, wire2832, wire2833, wire2834, wire2835, wire2836, wire2837, wire2838, wire2839, wire2840, wire2841, wire2842, wire2843, wire2844, wire2845, wire2846, wire2847, wire2848, wire2849, wire2850, wire2851, wire2852, wire2853, wire2854, wire2855, wire2856, wire2857, wire2858, wire2859, wire2860, wire2861, wire2862, wire2863, wire2864, wire2865, wire2866, wire2867, wire2868, wire2869, wire2870, wire2871, wire2872, wire2873, wire2874, wire2875, wire2876, wire2877, wire2878, wire2879, wire2880, wire2881, wire2882, wire2883, wire2884, wire2885, wire2886, wire2887, wire2888, wire2889, wire2890, wire2891, wire2892, wire2893, wire2894, wire2895, wire2896, wire2897, wire2898, wire2899, wire2900, wire2901, wire2902, wire2903, wire2904, wire2905, wire2906, wire2907, wire2908, wire2909, wire2910, wire2911, wire2912, wire2913, wire2914, wire2915, wire2916, wire2917, wire2918, wire2919, wire2920, wire2921, wire2922, wire2923, wire2924, wire2925, wire2926, wire2927, wire2928, wire2929, wire2930, wire2931, wire2932, wire2933, wire2934, wire2935, wire2936, wire2937, wire2938, wire2939, wire2940, wire2941, wire2942, wire2943, wire2944, wire2945, wire2946, wire2947, wire2948, wire2949, wire2950, wire2951, wire2952, wire2953, wire2954, wire2955, wire2956, wire2957, wire2958, wire2959, wire2960, wire2961, wire2962, wire2963, wire2964, wire2965, wire2966, wire2967, wire2968, wire2969, wire2970, wire2971, wire2972, wire2973, wire2974, wire2975, wire2976, wire2977, wire2978, wire2979, wire2980, wire2981, wire2982, wire2983, wire2984, wire2985, wire2986, wire2987, wire2988, wire2989, wire2990, wire2991, wire2992, wire2993, wire2994, wire2995, wire2996, wire2997, wire2998, wire2999, wire3000, wire3001, wire3002, wire3003, wire3004, wire3005, wire3006, wire3007, wire3008, wire3009, wire3010, wire3011, wire3012, wire3013, wire3014, wire3015, wire3016, wire3017, wire3018, wire3019, wire3020, wire3021, wire3022, wire3023, wire3024, wire3025, wire3026, wire3027, wire3028, wire3029, wire3030, wire3031, wire3032, wire3033, wire3034, wire3035, wire3036, wire3037, wire3038, wire3039, wire3040, wire3041, wire3042, wire3043, wire3044, wire3045, wire3046, wire3047, wire3048, wire3049, wire3050, wire3051, wire3052, wire3053, wire3054, wire3055, wire3056, wire3057, wire3058, wire3059, wire3060, wire3061, wire3062, wire3063, wire3064, wire3065, wire3066, wire3067, wire3068, wire3069, wire3070, wire3071, wire3072, wire3073, wire3074, wire3075, wire3076, wire3077, wire3078, wire3079, wire3080, wire3081, wire3082, wire3083, wire3084, wire3085, wire3086, wire3087, wire3088, wire3089, wire3090, wire3091, wire3092, wire3093, wire3094, wire3095, wire3096, wire3097, wire3098, wire3099, wire3100, wire3101, wire3102, wire3103, wire3104, wire3105, wire3106, wire3107, wire3108, wire3109, wire3110, wire3111, wire3112, wire3113, wire3114, wire3115, wire3116, wire3117, wire3118, wire3119, wire3120, wire3121, wire3122, wire3123, wire3124, wire3125, wire3126, wire3127, wire3128, wire3129, wire3130, wire3131, wire3132, wire3133, wire3134, wire3135, wire3136, wire3137, wire3138, wire3139, wire3140, wire3141, wire3142, wire3143, wire3144, wire3145, wire3146, wire3147, wire3148, wire3149, wire3150, wire3151, wire3152, wire3153, wire3154, wire3155, wire3156, wire3157, wire3158, wire3159, wire3160, wire3161, wire3162, wire3163, wire3164, wire3165, wire3166, wire3167, wire3168, wire3169, wire3170, wire3171, wire3172, wire3173, wire3174, wire3175, wire3176, wire3177, wire3178, wire3179, wire3180, wire3181, wire3182, wire3183, wire3184, wire3185, wire3186, wire3187, wire3188, wire3189, wire3190, wire3191, wire3192, wire3193, wire3194, wire3195, wire3196, wire3197, wire3198, wire3199, wire3200, wire3201, wire3202, wire3203, wire3204, wire3205, wire3206, wire3207, wire3208, wire3209, wire3210, wire3211, wire3212, wire3213, wire3214, wire3215, wire3216, wire3217, wire3218, wire3219, wire3220, wire3221, wire3222, wire3223, wire3224, wire3225, wire3226, wire3227, wire3228, wire3229, wire3230, wire3231, wire3232, wire3233, wire3234, wire3235, wire3236, wire3237, wire3238, wire3239, wire3240, wire3241, wire3242, wire3243, wire3244, wire3245, wire3246, wire3247, wire3248, wire3249, wire3250, wire3251, wire3252, wire3253, wire3254, wire3255, wire3256, wire3257, wire3258, wire3259, wire3260, wire3261, wire3262, wire3263, wire3264, wire3265, wire3266, wire3267, wire3268, wire3269, wire3270, wire3271, wire3272, wire3273, wire3274, wire3275, wire3276, wire3277, wire3278, wire3279, wire3280, wire3281, wire3282, wire3283, wire3284, wire3285, wire3286, wire3287, wire3288, wire3289, wire3290, wire3291, wire3292, wire3293, wire3294, wire3295, wire3296, wire3297, wire3298, wire3299, wire3300, wire3301, wire3302, wire3303, wire3304, wire3305, wire3306, wire3307, wire3308, wire3309, wire3310, wire3311, wire3312, wire3313, wire3314, wire3315, wire3316, wire3317, wire3318, wire3319, wire3320, wire3321, wire3322, wire3323, wire3324, wire3325, wire3326, wire3327, wire3328, wire3329, wire3330, wire3331, wire3332, wire3333, wire3334, wire3335, wire3336, wire3337, wire3338, wire3339, wire3340, wire3341, wire3342, wire3343, wire3344, wire3345, wire3346, wire3347, wire3348, wire3349, wire3350, wire3351, wire3352, wire3353, wire3354, wire3355, wire3356, wire3357, wire3358, wire3359, wire3360, wire3361, wire3362, wire3363, wire3364, wire3365, wire3366, wire3367, wire3368, wire3369, wire3370, wire3371, wire3372, wire3373, wire3374, wire3375, wire3376, wire3377, wire3378, wire3379, wire3380, wire3381, wire3382, wire3383, wire3384, wire3385, wire3386, wire3387, wire3388, wire3389, wire3390, wire3391, wire3392, wire3393, wire3394, wire3395, wire3396, wire3397, wire3398, wire3399, wire3400, wire3401, wire3402, wire3403, wire3404, wire3405, wire3406, wire3407, wire3408, wire3409, wire3410, wire3411, wire3412, wire3413, wire3414, wire3415, wire3416, wire3417, wire3418, wire3419, wire3420, wire3421, wire3422, wire3423, wire3424, wire3425, wire3426, wire3427, wire3428, wire3429, wire3430, wire3431, wire3432, wire3433, wire3434, wire3435, wire3436, wire3437, wire3438, wire3439, wire3440, wire3441, wire3442, wire3443, wire3444, wire3445, wire3446, wire3447, wire3448, wire3449, wire3450, wire3451, wire3452, wire3453, wire3454, wire3455, wire3456, wire3457, wire3458, wire3459, wire3460, wire3461, wire3462, wire3463, wire3464, wire3465, wire3466, wire3467, wire3468, wire3469, wire3470, wire3471, wire3472, wire3473, wire3474, wire3475, wire3476, wire3477, wire3478, wire3479, wire3480, wire3481, wire3482, wire3483, wire3484, wire3485, wire3486, wire3487, wire3488, wire3489, wire3490, wire3491, wire3492, wire3493, wire3494, wire3495, wire3496, wire3497, wire3498, wire3499, wire3500, wire3501, wire3502, wire3503, wire3504, wire3505, wire3506, wire3507, wire3508, wire3509, wire3510, wire3511, wire3512, wire3513, wire3514, wire3515, wire3516, wire3517, wire3518, wire3519, wire3520, wire3521, wire3522, wire3523, wire3524, wire3525, wire3526, wire3527, wire3528, wire3529, wire3530, wire3531, wire3532, wire3533, wire3534, wire3535, wire3536, wire3537, wire3538, wire3539, wire3540, wire3541, wire3542, wire3543, wire3544, wire3545, wire3546, wire3547, wire3548, wire3549, wire3550, wire3551, wire3552, wire3553, wire3554, wire3555, wire3556, wire3557, wire3558, wire3559, wire3560, wire3561, wire3562, wire3563, wire3564, wire3565, wire3566, wire3567, wire3568, wire3569, wire3570, wire3571, wire3572, wire3573, wire3574, wire3575, wire3576, wire3577, wire3578, wire3579, wire3580, wire3581, wire3582, wire3583, wire3584, wire3585, wire3586, wire3587, wire3588, wire3589, wire3590, wire3591, wire3592, wire3593, wire3594, wire3595, wire3596, wire3597, wire3598, wire3599, wire3600, wire3601, wire3602, wire3603, wire3604, wire3605, wire3606, wire3607, wire3608, wire3609, wire3610, wire3611, wire3612, wire3613, wire3614, wire3615, wire3616, wire3617, wire3618, wire3619, wire3620, wire3621, wire3622, wire3623, wire3624, wire3625, wire3626, wire3627, wire3628, wire3629, wire3630, wire3631, wire3632, wire3633, wire3634, wire3635, wire3636, wire3637, wire3638, wire3639, wire3640, wire3641, wire3642, wire3643, wire3644, wire3645, wire3646, wire3647, wire3648, wire3649, wire3650, wire3651, wire3652, wire3653, wire3654, wire3655, wire3656, wire3657, wire3658, wire3659, wire3660, wire3661, wire3662, wire3663, wire3664, wire3665, wire3666, wire3667, wire3668, wire3669, wire3670, wire3671, wire3672, wire3673, wire3674, wire3675, wire3676, wire3677, wire3678, wire3679, wire3680, wire3681, wire3682, wire3683, wire3684, wire3685, wire3686, wire3687, wire3688, wire3689, wire3690, wire3691, wire3692, wire3693, wire3694, wire3695, wire3696, wire3697, wire3698, wire3699, wire3700, wire3701, wire3702, wire3703, wire3704, wire3705, wire3706, wire3707, wire3708, wire3709, wire3710, wire3711, wire3712, wire3713, wire3714, wire3715, wire3716, wire3717, wire3718, wire3719, wire3720, wire3721, wire3722, wire3723, wire3724, wire3725, wire3726, wire3727, wire3728, wire3729, wire3730, wire3731, wire3732, wire3733, wire3734, wire3735, wire3736, wire3737, wire3738, wire3739, wire3740, wire3741, wire3742, wire3743, wire3744, wire3745, wire3746, wire3747, wire3748, wire3749, wire3750, wire3751, wire3752, wire3753, wire3754, wire3755, wire3756, wire3757, wire3758, wire3759, wire3760, wire3761, wire3762, wire3763, wire3764, wire3765, wire3766, wire3767, wire3768, wire3769, wire3770, wire3771, wire3772, wire3773, wire3774, wire3775, wire3776, wire3777, wire3778, wire3779, wire3780, wire3781, wire3782, wire3783, wire3784, wire3785, wire3786, wire3787, wire3788, wire3789, wire3790, wire3791, wire3792, wire3793, wire3794, wire3795, wire3796, wire3797, wire3798, wire3799, wire3800, wire3801, wire3802, wire3803, wire3804, wire3805, wire3806, wire3807, wire3808, wire3809, wire3810, wire3811, wire3812, wire3813, wire3814, wire3815, wire3816, wire3817, wire3818, wire3819, wire3820, wire3821, wire3822, wire3823, wire3824, wire3825, wire3826, wire3827, wire3828, wire3829, wire3830, wire3831, wire3832, wire3833, wire3834, wire3835, wire3836, wire3837, wire3838, wire3839, wire3840, wire3841, wire3842, wire3843, wire3844, wire3845, wire3846, wire3847, wire3848, wire3849, wire3850, wire3851, wire3852, wire3853, wire3854, wire3855, wire3856, wire3857, wire3858, wire3859, wire3860, wire3861, wire3862, wire3863, wire3864, wire3865, wire3866, wire3867, wire3868, wire3869, wire3870, wire3871, wire3872, wire3873, wire3874, wire3875, wire3876, wire3877, wire3878, wire3879, wire3880, wire3881, wire3882, wire3883, wire3884, wire3885, wire3886, wire3887, wire3888, wire3889, wire3890, wire3891, wire3892, wire3893, wire3894, wire3895, wire3896, wire3897, wire3898, wire3899, wire3900, wire3901, wire3902, wire3903, wire3904, wire3905, wire3906, wire3907, wire3908, wire3909, wire3910, wire3911, wire3912, wire3913, wire3914, wire3915, wire3916, wire3917, wire3918, wire3919, wire3920, wire3921, wire3922, wire3923, wire3924, wire3925, wire3926, wire3927, wire3928, wire3929, wire3930, wire3931, wire3932, wire3933, wire3934, wire3935, wire3936, wire3937, wire3938, wire3939, wire3940, wire3941, wire3942, wire3943, wire3944, wire3945, wire3946, wire3947, wire3948, wire3949, wire3950, wire3951, wire3952, wire3953, wire3954, wire3955, wire3956, wire3957, wire3958, wire3959, wire3960, wire3961, wire3962, wire3963, wire3964, wire3965, wire3966, wire3967, wire3968, wire3969, wire3970, wire3971, wire3972, wire3973, wire3974, wire3975, wire3976, wire3977, wire3978, wire3979, wire3980, wire3981, wire3982, wire3983, wire3984, wire3985, wire3986, wire3987, wire3988, wire3989, wire3990, wire3991, wire3992, wire3993, wire3994, wire3995, wire3996, wire3997, wire3998, wire3999, wire4000, wire4001, wire4002, wire4003, wire4004, wire4005, wire4006, wire4007, wire4008, wire4009, wire4010, wire4011, wire4012, wire4013, wire4014, wire4015, wire4016, wire4017, wire4018, wire4019, wire4020, wire4021, wire4022, wire4023, wire4024, wire4025, wire4026, wire4027, wire4028, wire4029, wire4030, wire4031, wire4032, wire4033, wire4034, wire4035, wire4036, wire4037, wire4038, wire4039, wire4040, wire4041, wire4042, wire4043, wire4044, wire4045, wire4046, wire4047, wire4048, wire4049, wire4050, wire4051, wire4052, wire4053, wire4054, wire4055, wire4056, wire4057, wire4058, wire4059, wire4060, wire4061, wire4062, wire4063, wire4064, wire4065, wire4066, wire4067, wire4068, wire4069, wire4070, wire4071, wire4072, wire4073, wire4074, wire4075, wire4076, wire4077, wire4078, wire4079, wire4080, wire4081, wire4082, wire4083, wire4084, wire4085, wire4086, wire4087, wire4088, wire4089, wire4090, wire4091, wire4092, wire4093, wire4094, wire4095;
    bufferH4096_12b$(.in(in), .out(buffered_input));
    assign wire0 = {4'd2, 4'd1};
    assign wire1 = {4'd2, 4'd1};
    assign wire2 = {4'd2, 4'd1};
    assign wire3 = {4'd2, 4'd1};
    assign wire4 = {4'd2, 4'd1};
    assign wire5 = {4'd2, 4'd1};
    assign wire6 = {4'd2, 4'd1};
    assign wire7 = {4'd2, 4'd1};
    assign wire8 = {4'd2, 4'd1};
    assign wire9 = {4'd2, 4'd1};
    assign wire10 = {4'd2, 4'd1};
    assign wire11 = {4'd2, 4'd1};
    assign wire12 = {4'd2, 4'd1};
    assign wire13 = {4'd2, 4'd1};
    assign wire14 = {4'd2, 4'd1};
    assign wire15 = {4'd2, 4'd1};
    assign wire16 = {4'd2, 4'd1};
    assign wire17 = {4'd2, 4'd1};
    assign wire18 = {4'd2, 4'd1};
    assign wire19 = {4'd2, 4'd1};
    assign wire20 = {4'd2, 4'd1};
    assign wire21 = {4'd2, 4'd1};
    assign wire22 = {4'd2, 4'd1};
    assign wire23 = {4'd2, 4'd1};
    assign wire24 = {4'd2, 4'd1};
    assign wire25 = {4'd2, 4'd1};
    assign wire26 = {4'd2, 4'd1};
    assign wire27 = {4'd2, 4'd1};
    assign wire28 = {4'd2, 4'd1};
    assign wire29 = {4'd2, 4'd1};
    assign wire30 = {4'd2, 4'd1};
    assign wire31 = {4'd2, 4'd1};
    assign wire32 = {4'd3, 4'd1};
    assign wire33 = {4'd3, 4'd1};
    assign wire34 = {4'd3, 4'd1};
    assign wire35 = {4'd3, 4'd1};
    assign wire36 = {4'd3, 4'd1};
    assign wire37 = {4'd3, 4'd1};
    assign wire38 = {4'd3, 4'd1};
    assign wire39 = {4'd3, 4'd1};
    assign wire40 = {4'd3, 4'd1};
    assign wire41 = {4'd3, 4'd1};
    assign wire42 = {4'd3, 4'd1};
    assign wire43 = {4'd3, 4'd1};
    assign wire44 = {4'd3, 4'd1};
    assign wire45 = {4'd3, 4'd1};
    assign wire46 = {4'd3, 4'd1};
    assign wire47 = {4'd3, 4'd1};
    assign wire48 = {4'd3, 4'd1};
    assign wire49 = {4'd3, 4'd1};
    assign wire50 = {4'd3, 4'd1};
    assign wire51 = {4'd3, 4'd1};
    assign wire52 = {4'd3, 4'd1};
    assign wire53 = {4'd3, 4'd1};
    assign wire54 = {4'd3, 4'd1};
    assign wire55 = {4'd3, 4'd1};
    assign wire56 = {4'd3, 4'd1};
    assign wire57 = {4'd3, 4'd1};
    assign wire58 = {4'd3, 4'd1};
    assign wire59 = {4'd3, 4'd1};
    assign wire60 = {4'd3, 4'd1};
    assign wire61 = {4'd3, 4'd1};
    assign wire62 = {4'd3, 4'd1};
    assign wire63 = {4'd3, 4'd1};
    assign wire64 = {4'd5, 4'd1};
    assign wire65 = {4'd5, 4'd1};
    assign wire66 = {4'd5, 4'd1};
    assign wire67 = {4'd5, 4'd1};
    assign wire68 = {4'd5, 4'd1};
    assign wire69 = {4'd5, 4'd1};
    assign wire70 = {4'd5, 4'd1};
    assign wire71 = {4'd5, 4'd1};
    assign wire72 = {4'd5, 4'd1};
    assign wire73 = {4'd5, 4'd1};
    assign wire74 = {4'd5, 4'd1};
    assign wire75 = {4'd5, 4'd1};
    assign wire76 = {4'd5, 4'd1};
    assign wire77 = {4'd5, 4'd1};
    assign wire78 = {4'd5, 4'd1};
    assign wire79 = {4'd5, 4'd1};
    assign wire80 = {4'd5, 4'd1};
    assign wire81 = {4'd5, 4'd1};
    assign wire82 = {4'd5, 4'd1};
    assign wire83 = {4'd5, 4'd1};
    assign wire84 = {4'd5, 4'd1};
    assign wire85 = {4'd5, 4'd1};
    assign wire86 = {4'd5, 4'd1};
    assign wire87 = {4'd5, 4'd1};
    assign wire88 = {4'd5, 4'd1};
    assign wire89 = {4'd5, 4'd1};
    assign wire90 = {4'd5, 4'd1};
    assign wire91 = {4'd5, 4'd1};
    assign wire92 = {4'd5, 4'd1};
    assign wire93 = {4'd5, 4'd1};
    assign wire94 = {4'd5, 4'd1};
    assign wire95 = {4'd5, 4'd1};
    assign wire96 = {4'd7, 4'd1};
    assign wire97 = {4'd7, 4'd1};
    assign wire98 = {4'd7, 4'd1};
    assign wire99 = {4'd7, 4'd1};
    assign wire100 = {4'd7, 4'd1};
    assign wire101 = {4'd7, 4'd1};
    assign wire102 = {4'd7, 4'd1};
    assign wire103 = {4'd7, 4'd1};
    assign wire104 = {4'd7, 4'd1};
    assign wire105 = {4'd7, 4'd1};
    assign wire106 = {4'd7, 4'd1};
    assign wire107 = {4'd7, 4'd1};
    assign wire108 = {4'd7, 4'd1};
    assign wire109 = {4'd7, 4'd1};
    assign wire110 = {4'd7, 4'd1};
    assign wire111 = {4'd7, 4'd1};
    assign wire112 = {4'd7, 4'd1};
    assign wire113 = {4'd7, 4'd1};
    assign wire114 = {4'd7, 4'd1};
    assign wire115 = {4'd7, 4'd1};
    assign wire116 = {4'd7, 4'd1};
    assign wire117 = {4'd7, 4'd1};
    assign wire118 = {4'd7, 4'd1};
    assign wire119 = {4'd7, 4'd1};
    assign wire120 = {4'd7, 4'd1};
    assign wire121 = {4'd7, 4'd1};
    assign wire122 = {4'd7, 4'd1};
    assign wire123 = {4'd7, 4'd1};
    assign wire124 = {4'd7, 4'd1};
    assign wire125 = {4'd7, 4'd1};
    assign wire126 = {4'd7, 4'd1};
    assign wire127 = {4'd7, 4'd1};
    assign wire128 = {4'd3, 4'd2};
    assign wire129 = {4'd3, 4'd2};
    assign wire130 = {4'd3, 4'd2};
    assign wire131 = {4'd3, 4'd2};
    assign wire132 = {4'd4, 4'd3};
    assign wire133 = {4'd7, 4'd6};
    assign wire134 = {4'd3, 4'd2};
    assign wire135 = {4'd3, 4'd2};
    assign wire136 = {4'd4, 4'd3};
    assign wire137 = {4'd4, 4'd3};
    assign wire138 = {4'd4, 4'd3};
    assign wire139 = {4'd4, 4'd3};
    assign wire140 = {4'd5, 4'd4};
    assign wire141 = {4'd4, 4'd3};
    assign wire142 = {4'd4, 4'd3};
    assign wire143 = {4'd4, 4'd3};
    assign wire144 = {4'd7, 4'd6};
    assign wire145 = {4'd7, 4'd6};
    assign wire146 = {4'd7, 4'd6};
    assign wire147 = {4'd7, 4'd6};
    assign wire148 = {4'd8, 4'd7};
    assign wire149 = {4'd7, 4'd6};
    assign wire150 = {4'd7, 4'd6};
    assign wire151 = {4'd7, 4'd6};
    assign wire152 = {4'd3, 4'd2};
    assign wire153 = {4'd3, 4'd2};
    assign wire154 = {4'd3, 4'd2};
    assign wire155 = {4'd3, 4'd2};
    assign wire156 = {4'd3, 4'd2};
    assign wire157 = {4'd3, 4'd2};
    assign wire158 = {4'd3, 4'd2};
    assign wire159 = {4'd3, 4'd2};
    assign wire160 = {4'd4, 4'd2};
    assign wire161 = {4'd4, 4'd2};
    assign wire162 = {4'd4, 4'd2};
    assign wire163 = {4'd4, 4'd2};
    assign wire164 = {4'd5, 4'd3};
    assign wire165 = {4'd8, 4'd6};
    assign wire166 = {4'd4, 4'd2};
    assign wire167 = {4'd4, 4'd2};
    assign wire168 = {4'd5, 4'd3};
    assign wire169 = {4'd5, 4'd3};
    assign wire170 = {4'd5, 4'd3};
    assign wire171 = {4'd5, 4'd3};
    assign wire172 = {4'd6, 4'd4};
    assign wire173 = {4'd5, 4'd3};
    assign wire174 = {4'd5, 4'd3};
    assign wire175 = {4'd5, 4'd3};
    assign wire176 = {4'd8, 4'd6};
    assign wire177 = {4'd8, 4'd6};
    assign wire178 = {4'd8, 4'd6};
    assign wire179 = {4'd8, 4'd6};
    assign wire180 = {4'd9, 4'd7};
    assign wire181 = {4'd8, 4'd6};
    assign wire182 = {4'd8, 4'd6};
    assign wire183 = {4'd8, 4'd6};
    assign wire184 = {4'd4, 4'd2};
    assign wire185 = {4'd4, 4'd2};
    assign wire186 = {4'd4, 4'd2};
    assign wire187 = {4'd4, 4'd2};
    assign wire188 = {4'd4, 4'd2};
    assign wire189 = {4'd4, 4'd2};
    assign wire190 = {4'd4, 4'd2};
    assign wire191 = {4'd4, 4'd2};
    assign wire192 = {4'd6, 4'd2};
    assign wire193 = {4'd6, 4'd2};
    assign wire194 = {4'd6, 4'd2};
    assign wire195 = {4'd6, 4'd2};
    assign wire196 = {4'd7, 4'd3};
    assign wire197 = {4'd10, 4'd6};
    assign wire198 = {4'd6, 4'd2};
    assign wire199 = {4'd6, 4'd2};
    assign wire200 = {4'd7, 4'd3};
    assign wire201 = {4'd7, 4'd3};
    assign wire202 = {4'd7, 4'd3};
    assign wire203 = {4'd7, 4'd3};
    assign wire204 = {4'd8, 4'd4};
    assign wire205 = {4'd7, 4'd3};
    assign wire206 = {4'd7, 4'd3};
    assign wire207 = {4'd7, 4'd3};
    assign wire208 = {4'd10, 4'd6};
    assign wire209 = {4'd10, 4'd6};
    assign wire210 = {4'd10, 4'd6};
    assign wire211 = {4'd10, 4'd6};
    assign wire212 = {4'd11, 4'd7};
    assign wire213 = {4'd10, 4'd6};
    assign wire214 = {4'd10, 4'd6};
    assign wire215 = {4'd10, 4'd6};
    assign wire216 = {4'd6, 4'd2};
    assign wire217 = {4'd6, 4'd2};
    assign wire218 = {4'd6, 4'd2};
    assign wire219 = {4'd6, 4'd2};
    assign wire220 = {4'd6, 4'd2};
    assign wire221 = {4'd6, 4'd2};
    assign wire222 = {4'd6, 4'd2};
    assign wire223 = {4'd6, 4'd2};
    assign wire224 = {4'd8, 4'd2};
    assign wire225 = {4'd8, 4'd2};
    assign wire226 = {4'd8, 4'd2};
    assign wire227 = {4'd8, 4'd2};
    assign wire228 = {4'd9, 4'd3};
    assign wire229 = {4'd12, 4'd6};
    assign wire230 = {4'd8, 4'd2};
    assign wire231 = {4'd8, 4'd2};
    assign wire232 = {4'd9, 4'd3};
    assign wire233 = {4'd9, 4'd3};
    assign wire234 = {4'd9, 4'd3};
    assign wire235 = {4'd9, 4'd3};
    assign wire236 = {4'd10, 4'd4};
    assign wire237 = {4'd9, 4'd3};
    assign wire238 = {4'd9, 4'd3};
    assign wire239 = {4'd9, 4'd3};
    assign wire240 = {4'd12, 4'd6};
    assign wire241 = {4'd12, 4'd6};
    assign wire242 = {4'd12, 4'd6};
    assign wire243 = {4'd12, 4'd6};
    assign wire244 = {4'd13, 4'd7};
    assign wire245 = {4'd12, 4'd6};
    assign wire246 = {4'd12, 4'd6};
    assign wire247 = {4'd12, 4'd6};
    assign wire248 = {4'd8, 4'd2};
    assign wire249 = {4'd8, 4'd2};
    assign wire250 = {4'd8, 4'd2};
    assign wire251 = {4'd8, 4'd2};
    assign wire252 = {4'd8, 4'd2};
    assign wire253 = {4'd8, 4'd2};
    assign wire254 = {4'd8, 4'd2};
    assign wire255 = {4'd8, 4'd2};
    assign wire256 = {4'd3, 4'd2};
    assign wire257 = {4'd3, 4'd2};
    assign wire258 = {4'd3, 4'd2};
    assign wire259 = {4'd3, 4'd2};
    assign wire260 = {4'd3, 4'd2};
    assign wire261 = {4'd3, 4'd2};
    assign wire262 = {4'd3, 4'd2};
    assign wire263 = {4'd3, 4'd2};
    assign wire264 = {4'd3, 4'd2};
    assign wire265 = {4'd3, 4'd2};
    assign wire266 = {4'd3, 4'd2};
    assign wire267 = {4'd3, 4'd2};
    assign wire268 = {4'd3, 4'd2};
    assign wire269 = {4'd3, 4'd2};
    assign wire270 = {4'd3, 4'd2};
    assign wire271 = {4'd3, 4'd2};
    assign wire272 = {4'd3, 4'd2};
    assign wire273 = {4'd3, 4'd2};
    assign wire274 = {4'd3, 4'd2};
    assign wire275 = {4'd3, 4'd2};
    assign wire276 = {4'd3, 4'd2};
    assign wire277 = {4'd3, 4'd2};
    assign wire278 = {4'd3, 4'd2};
    assign wire279 = {4'd3, 4'd2};
    assign wire280 = {4'd3, 4'd2};
    assign wire281 = {4'd3, 4'd2};
    assign wire282 = {4'd3, 4'd2};
    assign wire283 = {4'd3, 4'd2};
    assign wire284 = {4'd3, 4'd2};
    assign wire285 = {4'd3, 4'd2};
    assign wire286 = {4'd3, 4'd2};
    assign wire287 = {4'd3, 4'd2};
    assign wire288 = {4'd4, 4'd2};
    assign wire289 = {4'd4, 4'd2};
    assign wire290 = {4'd4, 4'd2};
    assign wire291 = {4'd4, 4'd2};
    assign wire292 = {4'd4, 4'd2};
    assign wire293 = {4'd4, 4'd2};
    assign wire294 = {4'd4, 4'd2};
    assign wire295 = {4'd4, 4'd2};
    assign wire296 = {4'd4, 4'd2};
    assign wire297 = {4'd4, 4'd2};
    assign wire298 = {4'd4, 4'd2};
    assign wire299 = {4'd4, 4'd2};
    assign wire300 = {4'd4, 4'd2};
    assign wire301 = {4'd4, 4'd2};
    assign wire302 = {4'd4, 4'd2};
    assign wire303 = {4'd4, 4'd2};
    assign wire304 = {4'd4, 4'd2};
    assign wire305 = {4'd4, 4'd2};
    assign wire306 = {4'd4, 4'd2};
    assign wire307 = {4'd4, 4'd2};
    assign wire308 = {4'd4, 4'd2};
    assign wire309 = {4'd4, 4'd2};
    assign wire310 = {4'd4, 4'd2};
    assign wire311 = {4'd4, 4'd2};
    assign wire312 = {4'd4, 4'd2};
    assign wire313 = {4'd4, 4'd2};
    assign wire314 = {4'd4, 4'd2};
    assign wire315 = {4'd4, 4'd2};
    assign wire316 = {4'd4, 4'd2};
    assign wire317 = {4'd4, 4'd2};
    assign wire318 = {4'd4, 4'd2};
    assign wire319 = {4'd4, 4'd2};
    assign wire320 = {4'd6, 4'd2};
    assign wire321 = {4'd6, 4'd2};
    assign wire322 = {4'd6, 4'd2};
    assign wire323 = {4'd6, 4'd2};
    assign wire324 = {4'd6, 4'd2};
    assign wire325 = {4'd6, 4'd2};
    assign wire326 = {4'd6, 4'd2};
    assign wire327 = {4'd6, 4'd2};
    assign wire328 = {4'd6, 4'd2};
    assign wire329 = {4'd6, 4'd2};
    assign wire330 = {4'd6, 4'd2};
    assign wire331 = {4'd6, 4'd2};
    assign wire332 = {4'd6, 4'd2};
    assign wire333 = {4'd6, 4'd2};
    assign wire334 = {4'd6, 4'd2};
    assign wire335 = {4'd6, 4'd2};
    assign wire336 = {4'd6, 4'd2};
    assign wire337 = {4'd6, 4'd2};
    assign wire338 = {4'd6, 4'd2};
    assign wire339 = {4'd6, 4'd2};
    assign wire340 = {4'd6, 4'd2};
    assign wire341 = {4'd6, 4'd2};
    assign wire342 = {4'd6, 4'd2};
    assign wire343 = {4'd6, 4'd2};
    assign wire344 = {4'd6, 4'd2};
    assign wire345 = {4'd6, 4'd2};
    assign wire346 = {4'd6, 4'd2};
    assign wire347 = {4'd6, 4'd2};
    assign wire348 = {4'd6, 4'd2};
    assign wire349 = {4'd6, 4'd2};
    assign wire350 = {4'd6, 4'd2};
    assign wire351 = {4'd6, 4'd2};
    assign wire352 = {4'd8, 4'd2};
    assign wire353 = {4'd8, 4'd2};
    assign wire354 = {4'd8, 4'd2};
    assign wire355 = {4'd8, 4'd2};
    assign wire356 = {4'd8, 4'd2};
    assign wire357 = {4'd8, 4'd2};
    assign wire358 = {4'd8, 4'd2};
    assign wire359 = {4'd8, 4'd2};
    assign wire360 = {4'd8, 4'd2};
    assign wire361 = {4'd8, 4'd2};
    assign wire362 = {4'd8, 4'd2};
    assign wire363 = {4'd8, 4'd2};
    assign wire364 = {4'd8, 4'd2};
    assign wire365 = {4'd8, 4'd2};
    assign wire366 = {4'd8, 4'd2};
    assign wire367 = {4'd8, 4'd2};
    assign wire368 = {4'd8, 4'd2};
    assign wire369 = {4'd8, 4'd2};
    assign wire370 = {4'd8, 4'd2};
    assign wire371 = {4'd8, 4'd2};
    assign wire372 = {4'd8, 4'd2};
    assign wire373 = {4'd8, 4'd2};
    assign wire374 = {4'd8, 4'd2};
    assign wire375 = {4'd8, 4'd2};
    assign wire376 = {4'd8, 4'd2};
    assign wire377 = {4'd8, 4'd2};
    assign wire378 = {4'd8, 4'd2};
    assign wire379 = {4'd8, 4'd2};
    assign wire380 = {4'd8, 4'd2};
    assign wire381 = {4'd8, 4'd2};
    assign wire382 = {4'd8, 4'd2};
    assign wire383 = {4'd8, 4'd2};
    assign wire384 = {4'd4, 4'd3};
    assign wire385 = {4'd4, 4'd3};
    assign wire386 = {4'd4, 4'd3};
    assign wire387 = {4'd4, 4'd3};
    assign wire388 = {4'd5, 4'd4};
    assign wire389 = {4'd8, 4'd7};
    assign wire390 = {4'd4, 4'd3};
    assign wire391 = {4'd4, 4'd3};
    assign wire392 = {4'd5, 4'd4};
    assign wire393 = {4'd5, 4'd4};
    assign wire394 = {4'd5, 4'd4};
    assign wire395 = {4'd5, 4'd4};
    assign wire396 = {4'd6, 4'd5};
    assign wire397 = {4'd5, 4'd4};
    assign wire398 = {4'd5, 4'd4};
    assign wire399 = {4'd5, 4'd4};
    assign wire400 = {4'd8, 4'd7};
    assign wire401 = {4'd8, 4'd7};
    assign wire402 = {4'd8, 4'd7};
    assign wire403 = {4'd8, 4'd7};
    assign wire404 = {4'd9, 4'd8};
    assign wire405 = {4'd8, 4'd7};
    assign wire406 = {4'd8, 4'd7};
    assign wire407 = {4'd8, 4'd7};
    assign wire408 = {4'd4, 4'd3};
    assign wire409 = {4'd4, 4'd3};
    assign wire410 = {4'd4, 4'd3};
    assign wire411 = {4'd4, 4'd3};
    assign wire412 = {4'd4, 4'd3};
    assign wire413 = {4'd4, 4'd3};
    assign wire414 = {4'd4, 4'd3};
    assign wire415 = {4'd4, 4'd3};
    assign wire416 = {4'd5, 4'd3};
    assign wire417 = {4'd5, 4'd3};
    assign wire418 = {4'd5, 4'd3};
    assign wire419 = {4'd5, 4'd3};
    assign wire420 = {4'd6, 4'd4};
    assign wire421 = {4'd9, 4'd7};
    assign wire422 = {4'd5, 4'd3};
    assign wire423 = {4'd5, 4'd3};
    assign wire424 = {4'd6, 4'd4};
    assign wire425 = {4'd6, 4'd4};
    assign wire426 = {4'd6, 4'd4};
    assign wire427 = {4'd6, 4'd4};
    assign wire428 = {4'd7, 4'd5};
    assign wire429 = {4'd6, 4'd4};
    assign wire430 = {4'd6, 4'd4};
    assign wire431 = {4'd6, 4'd4};
    assign wire432 = {4'd9, 4'd7};
    assign wire433 = {4'd9, 4'd7};
    assign wire434 = {4'd9, 4'd7};
    assign wire435 = {4'd9, 4'd7};
    assign wire436 = {4'd10, 4'd8};
    assign wire437 = {4'd9, 4'd7};
    assign wire438 = {4'd9, 4'd7};
    assign wire439 = {4'd9, 4'd7};
    assign wire440 = {4'd5, 4'd3};
    assign wire441 = {4'd5, 4'd3};
    assign wire442 = {4'd5, 4'd3};
    assign wire443 = {4'd5, 4'd3};
    assign wire444 = {4'd5, 4'd3};
    assign wire445 = {4'd5, 4'd3};
    assign wire446 = {4'd5, 4'd3};
    assign wire447 = {4'd5, 4'd3};
    assign wire448 = {4'd7, 4'd3};
    assign wire449 = {4'd7, 4'd3};
    assign wire450 = {4'd7, 4'd3};
    assign wire451 = {4'd7, 4'd3};
    assign wire452 = {4'd8, 4'd4};
    assign wire453 = {4'd11, 4'd7};
    assign wire454 = {4'd7, 4'd3};
    assign wire455 = {4'd7, 4'd3};
    assign wire456 = {4'd8, 4'd4};
    assign wire457 = {4'd8, 4'd4};
    assign wire458 = {4'd8, 4'd4};
    assign wire459 = {4'd8, 4'd4};
    assign wire460 = {4'd9, 4'd5};
    assign wire461 = {4'd8, 4'd4};
    assign wire462 = {4'd8, 4'd4};
    assign wire463 = {4'd8, 4'd4};
    assign wire464 = {4'd11, 4'd7};
    assign wire465 = {4'd11, 4'd7};
    assign wire466 = {4'd11, 4'd7};
    assign wire467 = {4'd11, 4'd7};
    assign wire468 = {4'd12, 4'd8};
    assign wire469 = {4'd11, 4'd7};
    assign wire470 = {4'd11, 4'd7};
    assign wire471 = {4'd11, 4'd7};
    assign wire472 = {4'd7, 4'd3};
    assign wire473 = {4'd7, 4'd3};
    assign wire474 = {4'd7, 4'd3};
    assign wire475 = {4'd7, 4'd3};
    assign wire476 = {4'd7, 4'd3};
    assign wire477 = {4'd7, 4'd3};
    assign wire478 = {4'd7, 4'd3};
    assign wire479 = {4'd7, 4'd3};
    assign wire480 = {4'd9, 4'd3};
    assign wire481 = {4'd9, 4'd3};
    assign wire482 = {4'd9, 4'd3};
    assign wire483 = {4'd9, 4'd3};
    assign wire484 = {4'd10, 4'd4};
    assign wire485 = {4'd13, 4'd7};
    assign wire486 = {4'd9, 4'd3};
    assign wire487 = {4'd9, 4'd3};
    assign wire488 = {4'd10, 4'd4};
    assign wire489 = {4'd10, 4'd4};
    assign wire490 = {4'd10, 4'd4};
    assign wire491 = {4'd10, 4'd4};
    assign wire492 = {4'd11, 4'd5};
    assign wire493 = {4'd10, 4'd4};
    assign wire494 = {4'd10, 4'd4};
    assign wire495 = {4'd10, 4'd4};
    assign wire496 = {4'd13, 4'd7};
    assign wire497 = {4'd13, 4'd7};
    assign wire498 = {4'd13, 4'd7};
    assign wire499 = {4'd13, 4'd7};
    assign wire500 = {4'd14, 4'd8};
    assign wire501 = {4'd13, 4'd7};
    assign wire502 = {4'd13, 4'd7};
    assign wire503 = {4'd13, 4'd7};
    assign wire504 = {4'd9, 4'd3};
    assign wire505 = {4'd9, 4'd3};
    assign wire506 = {4'd9, 4'd3};
    assign wire507 = {4'd9, 4'd3};
    assign wire508 = {4'd9, 4'd3};
    assign wire509 = {4'd9, 4'd3};
    assign wire510 = {4'd9, 4'd3};
    assign wire511 = {4'd9, 4'd3};
    assign wire512 = {4'd3, 4'd2};
    assign wire513 = {4'd3, 4'd2};
    assign wire514 = {4'd3, 4'd2};
    assign wire515 = {4'd3, 4'd2};
    assign wire516 = {4'd3, 4'd2};
    assign wire517 = {4'd3, 4'd2};
    assign wire518 = {4'd3, 4'd2};
    assign wire519 = {4'd3, 4'd2};
    assign wire520 = {4'd3, 4'd2};
    assign wire521 = {4'd3, 4'd2};
    assign wire522 = {4'd3, 4'd2};
    assign wire523 = {4'd3, 4'd2};
    assign wire524 = {4'd3, 4'd2};
    assign wire525 = {4'd3, 4'd2};
    assign wire526 = {4'd3, 4'd2};
    assign wire527 = {4'd3, 4'd2};
    assign wire528 = {4'd3, 4'd2};
    assign wire529 = {4'd3, 4'd2};
    assign wire530 = {4'd3, 4'd2};
    assign wire531 = {4'd3, 4'd2};
    assign wire532 = {4'd3, 4'd2};
    assign wire533 = {4'd3, 4'd2};
    assign wire534 = {4'd3, 4'd2};
    assign wire535 = {4'd3, 4'd2};
    assign wire536 = {4'd3, 4'd2};
    assign wire537 = {4'd3, 4'd2};
    assign wire538 = {4'd3, 4'd2};
    assign wire539 = {4'd3, 4'd2};
    assign wire540 = {4'd3, 4'd2};
    assign wire541 = {4'd3, 4'd2};
    assign wire542 = {4'd3, 4'd2};
    assign wire543 = {4'd3, 4'd2};
    assign wire544 = {4'd4, 4'd2};
    assign wire545 = {4'd4, 4'd2};
    assign wire546 = {4'd4, 4'd2};
    assign wire547 = {4'd4, 4'd2};
    assign wire548 = {4'd4, 4'd2};
    assign wire549 = {4'd4, 4'd2};
    assign wire550 = {4'd4, 4'd2};
    assign wire551 = {4'd4, 4'd2};
    assign wire552 = {4'd4, 4'd2};
    assign wire553 = {4'd4, 4'd2};
    assign wire554 = {4'd4, 4'd2};
    assign wire555 = {4'd4, 4'd2};
    assign wire556 = {4'd4, 4'd2};
    assign wire557 = {4'd4, 4'd2};
    assign wire558 = {4'd4, 4'd2};
    assign wire559 = {4'd4, 4'd2};
    assign wire560 = {4'd4, 4'd2};
    assign wire561 = {4'd4, 4'd2};
    assign wire562 = {4'd4, 4'd2};
    assign wire563 = {4'd4, 4'd2};
    assign wire564 = {4'd4, 4'd2};
    assign wire565 = {4'd4, 4'd2};
    assign wire566 = {4'd4, 4'd2};
    assign wire567 = {4'd4, 4'd2};
    assign wire568 = {4'd4, 4'd2};
    assign wire569 = {4'd4, 4'd2};
    assign wire570 = {4'd4, 4'd2};
    assign wire571 = {4'd4, 4'd2};
    assign wire572 = {4'd4, 4'd2};
    assign wire573 = {4'd4, 4'd2};
    assign wire574 = {4'd4, 4'd2};
    assign wire575 = {4'd4, 4'd2};
    assign wire576 = {4'd6, 4'd2};
    assign wire577 = {4'd6, 4'd2};
    assign wire578 = {4'd6, 4'd2};
    assign wire579 = {4'd6, 4'd2};
    assign wire580 = {4'd6, 4'd2};
    assign wire581 = {4'd6, 4'd2};
    assign wire582 = {4'd6, 4'd2};
    assign wire583 = {4'd6, 4'd2};
    assign wire584 = {4'd6, 4'd2};
    assign wire585 = {4'd6, 4'd2};
    assign wire586 = {4'd6, 4'd2};
    assign wire587 = {4'd6, 4'd2};
    assign wire588 = {4'd6, 4'd2};
    assign wire589 = {4'd6, 4'd2};
    assign wire590 = {4'd6, 4'd2};
    assign wire591 = {4'd6, 4'd2};
    assign wire592 = {4'd6, 4'd2};
    assign wire593 = {4'd6, 4'd2};
    assign wire594 = {4'd6, 4'd2};
    assign wire595 = {4'd6, 4'd2};
    assign wire596 = {4'd6, 4'd2};
    assign wire597 = {4'd6, 4'd2};
    assign wire598 = {4'd6, 4'd2};
    assign wire599 = {4'd6, 4'd2};
    assign wire600 = {4'd6, 4'd2};
    assign wire601 = {4'd6, 4'd2};
    assign wire602 = {4'd6, 4'd2};
    assign wire603 = {4'd6, 4'd2};
    assign wire604 = {4'd6, 4'd2};
    assign wire605 = {4'd6, 4'd2};
    assign wire606 = {4'd6, 4'd2};
    assign wire607 = {4'd6, 4'd2};
    assign wire608 = {4'd8, 4'd2};
    assign wire609 = {4'd8, 4'd2};
    assign wire610 = {4'd8, 4'd2};
    assign wire611 = {4'd8, 4'd2};
    assign wire612 = {4'd8, 4'd2};
    assign wire613 = {4'd8, 4'd2};
    assign wire614 = {4'd8, 4'd2};
    assign wire615 = {4'd8, 4'd2};
    assign wire616 = {4'd8, 4'd2};
    assign wire617 = {4'd8, 4'd2};
    assign wire618 = {4'd8, 4'd2};
    assign wire619 = {4'd8, 4'd2};
    assign wire620 = {4'd8, 4'd2};
    assign wire621 = {4'd8, 4'd2};
    assign wire622 = {4'd8, 4'd2};
    assign wire623 = {4'd8, 4'd2};
    assign wire624 = {4'd8, 4'd2};
    assign wire625 = {4'd8, 4'd2};
    assign wire626 = {4'd8, 4'd2};
    assign wire627 = {4'd8, 4'd2};
    assign wire628 = {4'd8, 4'd2};
    assign wire629 = {4'd8, 4'd2};
    assign wire630 = {4'd8, 4'd2};
    assign wire631 = {4'd8, 4'd2};
    assign wire632 = {4'd8, 4'd2};
    assign wire633 = {4'd8, 4'd2};
    assign wire634 = {4'd8, 4'd2};
    assign wire635 = {4'd8, 4'd2};
    assign wire636 = {4'd8, 4'd2};
    assign wire637 = {4'd8, 4'd2};
    assign wire638 = {4'd8, 4'd2};
    assign wire639 = {4'd8, 4'd2};
    assign wire640 = {4'd4, 4'd3};
    assign wire641 = {4'd4, 4'd3};
    assign wire642 = {4'd4, 4'd3};
    assign wire643 = {4'd4, 4'd3};
    assign wire644 = {4'd4, 4'd3};
    assign wire645 = {4'd6, 4'd5};
    assign wire646 = {4'd4, 4'd3};
    assign wire647 = {4'd4, 4'd3};
    assign wire648 = {4'd5, 4'd4};
    assign wire649 = {4'd5, 4'd4};
    assign wire650 = {4'd5, 4'd4};
    assign wire651 = {4'd5, 4'd4};
    assign wire652 = {4'd5, 4'd4};
    assign wire653 = {4'd5, 4'd4};
    assign wire654 = {4'd5, 4'd4};
    assign wire655 = {4'd5, 4'd4};
    assign wire656 = {4'd6, 4'd5};
    assign wire657 = {4'd6, 4'd5};
    assign wire658 = {4'd6, 4'd5};
    assign wire659 = {4'd6, 4'd5};
    assign wire660 = {4'd6, 4'd5};
    assign wire661 = {4'd6, 4'd5};
    assign wire662 = {4'd6, 4'd5};
    assign wire663 = {4'd6, 4'd5};
    assign wire664 = {4'd4, 4'd3};
    assign wire665 = {4'd4, 4'd3};
    assign wire666 = {4'd4, 4'd3};
    assign wire667 = {4'd4, 4'd3};
    assign wire668 = {4'd4, 4'd3};
    assign wire669 = {4'd4, 4'd3};
    assign wire670 = {4'd4, 4'd3};
    assign wire671 = {4'd4, 4'd3};
    assign wire672 = {4'd5, 4'd3};
    assign wire673 = {4'd5, 4'd3};
    assign wire674 = {4'd5, 4'd3};
    assign wire675 = {4'd5, 4'd3};
    assign wire676 = {4'd5, 4'd3};
    assign wire677 = {4'd7, 4'd5};
    assign wire678 = {4'd5, 4'd3};
    assign wire679 = {4'd5, 4'd3};
    assign wire680 = {4'd6, 4'd4};
    assign wire681 = {4'd6, 4'd4};
    assign wire682 = {4'd6, 4'd4};
    assign wire683 = {4'd6, 4'd4};
    assign wire684 = {4'd6, 4'd4};
    assign wire685 = {4'd6, 4'd4};
    assign wire686 = {4'd6, 4'd4};
    assign wire687 = {4'd6, 4'd4};
    assign wire688 = {4'd7, 4'd5};
    assign wire689 = {4'd7, 4'd5};
    assign wire690 = {4'd7, 4'd5};
    assign wire691 = {4'd7, 4'd5};
    assign wire692 = {4'd7, 4'd5};
    assign wire693 = {4'd7, 4'd5};
    assign wire694 = {4'd7, 4'd5};
    assign wire695 = {4'd7, 4'd5};
    assign wire696 = {4'd5, 4'd3};
    assign wire697 = {4'd5, 4'd3};
    assign wire698 = {4'd5, 4'd3};
    assign wire699 = {4'd5, 4'd3};
    assign wire700 = {4'd5, 4'd3};
    assign wire701 = {4'd5, 4'd3};
    assign wire702 = {4'd5, 4'd3};
    assign wire703 = {4'd5, 4'd3};
    assign wire704 = {4'd7, 4'd3};
    assign wire705 = {4'd7, 4'd3};
    assign wire706 = {4'd7, 4'd3};
    assign wire707 = {4'd7, 4'd3};
    assign wire708 = {4'd7, 4'd3};
    assign wire709 = {4'd9, 4'd5};
    assign wire710 = {4'd7, 4'd3};
    assign wire711 = {4'd7, 4'd3};
    assign wire712 = {4'd8, 4'd4};
    assign wire713 = {4'd8, 4'd4};
    assign wire714 = {4'd8, 4'd4};
    assign wire715 = {4'd8, 4'd4};
    assign wire716 = {4'd8, 4'd4};
    assign wire717 = {4'd8, 4'd4};
    assign wire718 = {4'd8, 4'd4};
    assign wire719 = {4'd8, 4'd4};
    assign wire720 = {4'd9, 4'd5};
    assign wire721 = {4'd9, 4'd5};
    assign wire722 = {4'd9, 4'd5};
    assign wire723 = {4'd9, 4'd5};
    assign wire724 = {4'd9, 4'd5};
    assign wire725 = {4'd9, 4'd5};
    assign wire726 = {4'd9, 4'd5};
    assign wire727 = {4'd9, 4'd5};
    assign wire728 = {4'd7, 4'd3};
    assign wire729 = {4'd7, 4'd3};
    assign wire730 = {4'd7, 4'd3};
    assign wire731 = {4'd7, 4'd3};
    assign wire732 = {4'd7, 4'd3};
    assign wire733 = {4'd7, 4'd3};
    assign wire734 = {4'd7, 4'd3};
    assign wire735 = {4'd7, 4'd3};
    assign wire736 = {4'd9, 4'd3};
    assign wire737 = {4'd9, 4'd3};
    assign wire738 = {4'd9, 4'd3};
    assign wire739 = {4'd9, 4'd3};
    assign wire740 = {4'd9, 4'd3};
    assign wire741 = {4'd11, 4'd5};
    assign wire742 = {4'd9, 4'd3};
    assign wire743 = {4'd9, 4'd3};
    assign wire744 = {4'd10, 4'd4};
    assign wire745 = {4'd10, 4'd4};
    assign wire746 = {4'd10, 4'd4};
    assign wire747 = {4'd10, 4'd4};
    assign wire748 = {4'd10, 4'd4};
    assign wire749 = {4'd10, 4'd4};
    assign wire750 = {4'd10, 4'd4};
    assign wire751 = {4'd10, 4'd4};
    assign wire752 = {4'd11, 4'd5};
    assign wire753 = {4'd11, 4'd5};
    assign wire754 = {4'd11, 4'd5};
    assign wire755 = {4'd11, 4'd5};
    assign wire756 = {4'd11, 4'd5};
    assign wire757 = {4'd11, 4'd5};
    assign wire758 = {4'd11, 4'd5};
    assign wire759 = {4'd11, 4'd5};
    assign wire760 = {4'd9, 4'd3};
    assign wire761 = {4'd9, 4'd3};
    assign wire762 = {4'd9, 4'd3};
    assign wire763 = {4'd9, 4'd3};
    assign wire764 = {4'd9, 4'd3};
    assign wire765 = {4'd9, 4'd3};
    assign wire766 = {4'd9, 4'd3};
    assign wire767 = {4'd9, 4'd3};
    assign wire768 = {4'd4, 4'd3};
    assign wire769 = {4'd4, 4'd3};
    assign wire770 = {4'd4, 4'd3};
    assign wire771 = {4'd4, 4'd3};
    assign wire772 = {4'd4, 4'd3};
    assign wire773 = {4'd4, 4'd3};
    assign wire774 = {4'd4, 4'd3};
    assign wire775 = {4'd4, 4'd3};
    assign wire776 = {4'd4, 4'd3};
    assign wire777 = {4'd4, 4'd3};
    assign wire778 = {4'd4, 4'd3};
    assign wire779 = {4'd4, 4'd3};
    assign wire780 = {4'd4, 4'd3};
    assign wire781 = {4'd4, 4'd3};
    assign wire782 = {4'd4, 4'd3};
    assign wire783 = {4'd4, 4'd3};
    assign wire784 = {4'd4, 4'd3};
    assign wire785 = {4'd4, 4'd3};
    assign wire786 = {4'd4, 4'd3};
    assign wire787 = {4'd4, 4'd3};
    assign wire788 = {4'd4, 4'd3};
    assign wire789 = {4'd4, 4'd3};
    assign wire790 = {4'd4, 4'd3};
    assign wire791 = {4'd4, 4'd3};
    assign wire792 = {4'd4, 4'd3};
    assign wire793 = {4'd4, 4'd3};
    assign wire794 = {4'd4, 4'd3};
    assign wire795 = {4'd4, 4'd3};
    assign wire796 = {4'd4, 4'd3};
    assign wire797 = {4'd4, 4'd3};
    assign wire798 = {4'd4, 4'd3};
    assign wire799 = {4'd4, 4'd3};
    assign wire800 = {4'd5, 4'd3};
    assign wire801 = {4'd5, 4'd3};
    assign wire802 = {4'd5, 4'd3};
    assign wire803 = {4'd5, 4'd3};
    assign wire804 = {4'd5, 4'd3};
    assign wire805 = {4'd5, 4'd3};
    assign wire806 = {4'd5, 4'd3};
    assign wire807 = {4'd5, 4'd3};
    assign wire808 = {4'd5, 4'd3};
    assign wire809 = {4'd5, 4'd3};
    assign wire810 = {4'd5, 4'd3};
    assign wire811 = {4'd5, 4'd3};
    assign wire812 = {4'd5, 4'd3};
    assign wire813 = {4'd5, 4'd3};
    assign wire814 = {4'd5, 4'd3};
    assign wire815 = {4'd5, 4'd3};
    assign wire816 = {4'd5, 4'd3};
    assign wire817 = {4'd5, 4'd3};
    assign wire818 = {4'd5, 4'd3};
    assign wire819 = {4'd5, 4'd3};
    assign wire820 = {4'd5, 4'd3};
    assign wire821 = {4'd5, 4'd3};
    assign wire822 = {4'd5, 4'd3};
    assign wire823 = {4'd5, 4'd3};
    assign wire824 = {4'd5, 4'd3};
    assign wire825 = {4'd5, 4'd3};
    assign wire826 = {4'd5, 4'd3};
    assign wire827 = {4'd5, 4'd3};
    assign wire828 = {4'd5, 4'd3};
    assign wire829 = {4'd5, 4'd3};
    assign wire830 = {4'd5, 4'd3};
    assign wire831 = {4'd5, 4'd3};
    assign wire832 = {4'd7, 4'd3};
    assign wire833 = {4'd7, 4'd3};
    assign wire834 = {4'd7, 4'd3};
    assign wire835 = {4'd7, 4'd3};
    assign wire836 = {4'd7, 4'd3};
    assign wire837 = {4'd7, 4'd3};
    assign wire838 = {4'd7, 4'd3};
    assign wire839 = {4'd7, 4'd3};
    assign wire840 = {4'd7, 4'd3};
    assign wire841 = {4'd7, 4'd3};
    assign wire842 = {4'd7, 4'd3};
    assign wire843 = {4'd7, 4'd3};
    assign wire844 = {4'd7, 4'd3};
    assign wire845 = {4'd7, 4'd3};
    assign wire846 = {4'd7, 4'd3};
    assign wire847 = {4'd7, 4'd3};
    assign wire848 = {4'd7, 4'd3};
    assign wire849 = {4'd7, 4'd3};
    assign wire850 = {4'd7, 4'd3};
    assign wire851 = {4'd7, 4'd3};
    assign wire852 = {4'd7, 4'd3};
    assign wire853 = {4'd7, 4'd3};
    assign wire854 = {4'd7, 4'd3};
    assign wire855 = {4'd7, 4'd3};
    assign wire856 = {4'd7, 4'd3};
    assign wire857 = {4'd7, 4'd3};
    assign wire858 = {4'd7, 4'd3};
    assign wire859 = {4'd7, 4'd3};
    assign wire860 = {4'd7, 4'd3};
    assign wire861 = {4'd7, 4'd3};
    assign wire862 = {4'd7, 4'd3};
    assign wire863 = {4'd7, 4'd3};
    assign wire864 = {4'd9, 4'd3};
    assign wire865 = {4'd9, 4'd3};
    assign wire866 = {4'd9, 4'd3};
    assign wire867 = {4'd9, 4'd3};
    assign wire868 = {4'd9, 4'd3};
    assign wire869 = {4'd9, 4'd3};
    assign wire870 = {4'd9, 4'd3};
    assign wire871 = {4'd9, 4'd3};
    assign wire872 = {4'd9, 4'd3};
    assign wire873 = {4'd9, 4'd3};
    assign wire874 = {4'd9, 4'd3};
    assign wire875 = {4'd9, 4'd3};
    assign wire876 = {4'd9, 4'd3};
    assign wire877 = {4'd9, 4'd3};
    assign wire878 = {4'd9, 4'd3};
    assign wire879 = {4'd9, 4'd3};
    assign wire880 = {4'd9, 4'd3};
    assign wire881 = {4'd9, 4'd3};
    assign wire882 = {4'd9, 4'd3};
    assign wire883 = {4'd9, 4'd3};
    assign wire884 = {4'd9, 4'd3};
    assign wire885 = {4'd9, 4'd3};
    assign wire886 = {4'd9, 4'd3};
    assign wire887 = {4'd9, 4'd3};
    assign wire888 = {4'd9, 4'd3};
    assign wire889 = {4'd9, 4'd3};
    assign wire890 = {4'd9, 4'd3};
    assign wire891 = {4'd9, 4'd3};
    assign wire892 = {4'd9, 4'd3};
    assign wire893 = {4'd9, 4'd3};
    assign wire894 = {4'd9, 4'd3};
    assign wire895 = {4'd9, 4'd3};
    assign wire896 = {4'd5, 4'd4};
    assign wire897 = {4'd5, 4'd4};
    assign wire898 = {4'd5, 4'd4};
    assign wire899 = {4'd5, 4'd4};
    assign wire900 = {4'd5, 4'd4};
    assign wire901 = {4'd7, 4'd6};
    assign wire902 = {4'd5, 4'd4};
    assign wire903 = {4'd5, 4'd4};
    assign wire904 = {4'd6, 4'd5};
    assign wire905 = {4'd6, 4'd5};
    assign wire906 = {4'd6, 4'd5};
    assign wire907 = {4'd6, 4'd5};
    assign wire908 = {4'd6, 4'd5};
    assign wire909 = {4'd6, 4'd5};
    assign wire910 = {4'd6, 4'd5};
    assign wire911 = {4'd6, 4'd5};
    assign wire912 = {4'd7, 4'd6};
    assign wire913 = {4'd7, 4'd6};
    assign wire914 = {4'd7, 4'd6};
    assign wire915 = {4'd7, 4'd6};
    assign wire916 = {4'd7, 4'd6};
    assign wire917 = {4'd7, 4'd6};
    assign wire918 = {4'd7, 4'd6};
    assign wire919 = {4'd7, 4'd6};
    assign wire920 = {4'd5, 4'd4};
    assign wire921 = {4'd5, 4'd4};
    assign wire922 = {4'd5, 4'd4};
    assign wire923 = {4'd5, 4'd4};
    assign wire924 = {4'd5, 4'd4};
    assign wire925 = {4'd5, 4'd4};
    assign wire926 = {4'd5, 4'd4};
    assign wire927 = {4'd5, 4'd4};
    assign wire928 = {4'd6, 4'd4};
    assign wire929 = {4'd6, 4'd4};
    assign wire930 = {4'd6, 4'd4};
    assign wire931 = {4'd6, 4'd4};
    assign wire932 = {4'd6, 4'd4};
    assign wire933 = {4'd8, 4'd6};
    assign wire934 = {4'd6, 4'd4};
    assign wire935 = {4'd6, 4'd4};
    assign wire936 = {4'd7, 4'd5};
    assign wire937 = {4'd7, 4'd5};
    assign wire938 = {4'd7, 4'd5};
    assign wire939 = {4'd7, 4'd5};
    assign wire940 = {4'd7, 4'd5};
    assign wire941 = {4'd7, 4'd5};
    assign wire942 = {4'd7, 4'd5};
    assign wire943 = {4'd7, 4'd5};
    assign wire944 = {4'd8, 4'd6};
    assign wire945 = {4'd8, 4'd6};
    assign wire946 = {4'd8, 4'd6};
    assign wire947 = {4'd8, 4'd6};
    assign wire948 = {4'd8, 4'd6};
    assign wire949 = {4'd8, 4'd6};
    assign wire950 = {4'd8, 4'd6};
    assign wire951 = {4'd8, 4'd6};
    assign wire952 = {4'd6, 4'd4};
    assign wire953 = {4'd6, 4'd4};
    assign wire954 = {4'd6, 4'd4};
    assign wire955 = {4'd6, 4'd4};
    assign wire956 = {4'd6, 4'd4};
    assign wire957 = {4'd6, 4'd4};
    assign wire958 = {4'd6, 4'd4};
    assign wire959 = {4'd6, 4'd4};
    assign wire960 = {4'd8, 4'd4};
    assign wire961 = {4'd8, 4'd4};
    assign wire962 = {4'd8, 4'd4};
    assign wire963 = {4'd8, 4'd4};
    assign wire964 = {4'd8, 4'd4};
    assign wire965 = {4'd10, 4'd6};
    assign wire966 = {4'd8, 4'd4};
    assign wire967 = {4'd8, 4'd4};
    assign wire968 = {4'd9, 4'd5};
    assign wire969 = {4'd9, 4'd5};
    assign wire970 = {4'd9, 4'd5};
    assign wire971 = {4'd9, 4'd5};
    assign wire972 = {4'd9, 4'd5};
    assign wire973 = {4'd9, 4'd5};
    assign wire974 = {4'd9, 4'd5};
    assign wire975 = {4'd9, 4'd5};
    assign wire976 = {4'd10, 4'd6};
    assign wire977 = {4'd10, 4'd6};
    assign wire978 = {4'd10, 4'd6};
    assign wire979 = {4'd10, 4'd6};
    assign wire980 = {4'd10, 4'd6};
    assign wire981 = {4'd10, 4'd6};
    assign wire982 = {4'd10, 4'd6};
    assign wire983 = {4'd10, 4'd6};
    assign wire984 = {4'd8, 4'd4};
    assign wire985 = {4'd8, 4'd4};
    assign wire986 = {4'd8, 4'd4};
    assign wire987 = {4'd8, 4'd4};
    assign wire988 = {4'd8, 4'd4};
    assign wire989 = {4'd8, 4'd4};
    assign wire990 = {4'd8, 4'd4};
    assign wire991 = {4'd8, 4'd4};
    assign wire992 = {4'd10, 4'd4};
    assign wire993 = {4'd10, 4'd4};
    assign wire994 = {4'd10, 4'd4};
    assign wire995 = {4'd10, 4'd4};
    assign wire996 = {4'd10, 4'd4};
    assign wire997 = {4'd12, 4'd6};
    assign wire998 = {4'd10, 4'd4};
    assign wire999 = {4'd10, 4'd4};
    assign wire1000 = {4'd11, 4'd5};
    assign wire1001 = {4'd11, 4'd5};
    assign wire1002 = {4'd11, 4'd5};
    assign wire1003 = {4'd11, 4'd5};
    assign wire1004 = {4'd11, 4'd5};
    assign wire1005 = {4'd11, 4'd5};
    assign wire1006 = {4'd11, 4'd5};
    assign wire1007 = {4'd11, 4'd5};
    assign wire1008 = {4'd12, 4'd6};
    assign wire1009 = {4'd12, 4'd6};
    assign wire1010 = {4'd12, 4'd6};
    assign wire1011 = {4'd12, 4'd6};
    assign wire1012 = {4'd12, 4'd6};
    assign wire1013 = {4'd12, 4'd6};
    assign wire1014 = {4'd12, 4'd6};
    assign wire1015 = {4'd12, 4'd6};
    assign wire1016 = {4'd10, 4'd4};
    assign wire1017 = {4'd10, 4'd4};
    assign wire1018 = {4'd10, 4'd4};
    assign wire1019 = {4'd10, 4'd4};
    assign wire1020 = {4'd10, 4'd4};
    assign wire1021 = {4'd10, 4'd4};
    assign wire1022 = {4'd10, 4'd4};
    assign wire1023 = {4'd10, 4'd4};
    assign wire1024 = {4'd3, 4'd2};
    assign wire1025 = {4'd3, 4'd2};
    assign wire1026 = {4'd3, 4'd2};
    assign wire1027 = {4'd3, 4'd2};
    assign wire1028 = {4'd3, 4'd2};
    assign wire1029 = {4'd3, 4'd2};
    assign wire1030 = {4'd3, 4'd2};
    assign wire1031 = {4'd3, 4'd2};
    assign wire1032 = {4'd3, 4'd2};
    assign wire1033 = {4'd3, 4'd2};
    assign wire1034 = {4'd3, 4'd2};
    assign wire1035 = {4'd3, 4'd2};
    assign wire1036 = {4'd3, 4'd2};
    assign wire1037 = {4'd3, 4'd2};
    assign wire1038 = {4'd3, 4'd2};
    assign wire1039 = {4'd3, 4'd2};
    assign wire1040 = {4'd3, 4'd2};
    assign wire1041 = {4'd3, 4'd2};
    assign wire1042 = {4'd3, 4'd2};
    assign wire1043 = {4'd3, 4'd2};
    assign wire1044 = {4'd3, 4'd2};
    assign wire1045 = {4'd3, 4'd2};
    assign wire1046 = {4'd3, 4'd2};
    assign wire1047 = {4'd3, 4'd2};
    assign wire1048 = {4'd3, 4'd2};
    assign wire1049 = {4'd3, 4'd2};
    assign wire1050 = {4'd3, 4'd2};
    assign wire1051 = {4'd3, 4'd2};
    assign wire1052 = {4'd3, 4'd2};
    assign wire1053 = {4'd3, 4'd2};
    assign wire1054 = {4'd3, 4'd2};
    assign wire1055 = {4'd3, 4'd2};
    assign wire1056 = {4'd4, 4'd2};
    assign wire1057 = {4'd4, 4'd2};
    assign wire1058 = {4'd4, 4'd2};
    assign wire1059 = {4'd4, 4'd2};
    assign wire1060 = {4'd4, 4'd2};
    assign wire1061 = {4'd4, 4'd2};
    assign wire1062 = {4'd4, 4'd2};
    assign wire1063 = {4'd4, 4'd2};
    assign wire1064 = {4'd4, 4'd2};
    assign wire1065 = {4'd4, 4'd2};
    assign wire1066 = {4'd4, 4'd2};
    assign wire1067 = {4'd4, 4'd2};
    assign wire1068 = {4'd4, 4'd2};
    assign wire1069 = {4'd4, 4'd2};
    assign wire1070 = {4'd4, 4'd2};
    assign wire1071 = {4'd4, 4'd2};
    assign wire1072 = {4'd4, 4'd2};
    assign wire1073 = {4'd4, 4'd2};
    assign wire1074 = {4'd4, 4'd2};
    assign wire1075 = {4'd4, 4'd2};
    assign wire1076 = {4'd4, 4'd2};
    assign wire1077 = {4'd4, 4'd2};
    assign wire1078 = {4'd4, 4'd2};
    assign wire1079 = {4'd4, 4'd2};
    assign wire1080 = {4'd4, 4'd2};
    assign wire1081 = {4'd4, 4'd2};
    assign wire1082 = {4'd4, 4'd2};
    assign wire1083 = {4'd4, 4'd2};
    assign wire1084 = {4'd4, 4'd2};
    assign wire1085 = {4'd4, 4'd2};
    assign wire1086 = {4'd4, 4'd2};
    assign wire1087 = {4'd4, 4'd2};
    assign wire1088 = {4'd6, 4'd2};
    assign wire1089 = {4'd6, 4'd2};
    assign wire1090 = {4'd6, 4'd2};
    assign wire1091 = {4'd6, 4'd2};
    assign wire1092 = {4'd6, 4'd2};
    assign wire1093 = {4'd6, 4'd2};
    assign wire1094 = {4'd6, 4'd2};
    assign wire1095 = {4'd6, 4'd2};
    assign wire1096 = {4'd6, 4'd2};
    assign wire1097 = {4'd6, 4'd2};
    assign wire1098 = {4'd6, 4'd2};
    assign wire1099 = {4'd6, 4'd2};
    assign wire1100 = {4'd6, 4'd2};
    assign wire1101 = {4'd6, 4'd2};
    assign wire1102 = {4'd6, 4'd2};
    assign wire1103 = {4'd6, 4'd2};
    assign wire1104 = {4'd6, 4'd2};
    assign wire1105 = {4'd6, 4'd2};
    assign wire1106 = {4'd6, 4'd2};
    assign wire1107 = {4'd6, 4'd2};
    assign wire1108 = {4'd6, 4'd2};
    assign wire1109 = {4'd6, 4'd2};
    assign wire1110 = {4'd6, 4'd2};
    assign wire1111 = {4'd6, 4'd2};
    assign wire1112 = {4'd6, 4'd2};
    assign wire1113 = {4'd6, 4'd2};
    assign wire1114 = {4'd6, 4'd2};
    assign wire1115 = {4'd6, 4'd2};
    assign wire1116 = {4'd6, 4'd2};
    assign wire1117 = {4'd6, 4'd2};
    assign wire1118 = {4'd6, 4'd2};
    assign wire1119 = {4'd6, 4'd2};
    assign wire1120 = {4'd8, 4'd2};
    assign wire1121 = {4'd8, 4'd2};
    assign wire1122 = {4'd8, 4'd2};
    assign wire1123 = {4'd8, 4'd2};
    assign wire1124 = {4'd8, 4'd2};
    assign wire1125 = {4'd8, 4'd2};
    assign wire1126 = {4'd8, 4'd2};
    assign wire1127 = {4'd8, 4'd2};
    assign wire1128 = {4'd8, 4'd2};
    assign wire1129 = {4'd8, 4'd2};
    assign wire1130 = {4'd8, 4'd2};
    assign wire1131 = {4'd8, 4'd2};
    assign wire1132 = {4'd8, 4'd2};
    assign wire1133 = {4'd8, 4'd2};
    assign wire1134 = {4'd8, 4'd2};
    assign wire1135 = {4'd8, 4'd2};
    assign wire1136 = {4'd8, 4'd2};
    assign wire1137 = {4'd8, 4'd2};
    assign wire1138 = {4'd8, 4'd2};
    assign wire1139 = {4'd8, 4'd2};
    assign wire1140 = {4'd8, 4'd2};
    assign wire1141 = {4'd8, 4'd2};
    assign wire1142 = {4'd8, 4'd2};
    assign wire1143 = {4'd8, 4'd2};
    assign wire1144 = {4'd8, 4'd2};
    assign wire1145 = {4'd8, 4'd2};
    assign wire1146 = {4'd8, 4'd2};
    assign wire1147 = {4'd8, 4'd2};
    assign wire1148 = {4'd8, 4'd2};
    assign wire1149 = {4'd8, 4'd2};
    assign wire1150 = {4'd8, 4'd2};
    assign wire1151 = {4'd8, 4'd2};
    assign wire1152 = {4'd4, 4'd3};
    assign wire1153 = {4'd4, 4'd3};
    assign wire1154 = {4'd4, 4'd3};
    assign wire1155 = {4'd4, 4'd3};
    assign wire1156 = {4'd5, 4'd4};
    assign wire1157 = {4'd8, 4'd7};
    assign wire1158 = {4'd4, 4'd3};
    assign wire1159 = {4'd4, 4'd3};
    assign wire1160 = {4'd5, 4'd4};
    assign wire1161 = {4'd5, 4'd4};
    assign wire1162 = {4'd5, 4'd4};
    assign wire1163 = {4'd5, 4'd4};
    assign wire1164 = {4'd6, 4'd5};
    assign wire1165 = {4'd5, 4'd4};
    assign wire1166 = {4'd5, 4'd4};
    assign wire1167 = {4'd5, 4'd4};
    assign wire1168 = {4'd8, 4'd7};
    assign wire1169 = {4'd8, 4'd7};
    assign wire1170 = {4'd8, 4'd7};
    assign wire1171 = {4'd8, 4'd7};
    assign wire1172 = {4'd9, 4'd8};
    assign wire1173 = {4'd8, 4'd7};
    assign wire1174 = {4'd8, 4'd7};
    assign wire1175 = {4'd8, 4'd7};
    assign wire1176 = {4'd4, 4'd3};
    assign wire1177 = {4'd4, 4'd3};
    assign wire1178 = {4'd4, 4'd3};
    assign wire1179 = {4'd4, 4'd3};
    assign wire1180 = {4'd4, 4'd3};
    assign wire1181 = {4'd4, 4'd3};
    assign wire1182 = {4'd4, 4'd3};
    assign wire1183 = {4'd4, 4'd3};
    assign wire1184 = {4'd5, 4'd3};
    assign wire1185 = {4'd5, 4'd3};
    assign wire1186 = {4'd5, 4'd3};
    assign wire1187 = {4'd5, 4'd3};
    assign wire1188 = {4'd6, 4'd4};
    assign wire1189 = {4'd9, 4'd7};
    assign wire1190 = {4'd5, 4'd3};
    assign wire1191 = {4'd5, 4'd3};
    assign wire1192 = {4'd6, 4'd4};
    assign wire1193 = {4'd6, 4'd4};
    assign wire1194 = {4'd6, 4'd4};
    assign wire1195 = {4'd6, 4'd4};
    assign wire1196 = {4'd7, 4'd5};
    assign wire1197 = {4'd6, 4'd4};
    assign wire1198 = {4'd6, 4'd4};
    assign wire1199 = {4'd6, 4'd4};
    assign wire1200 = {4'd9, 4'd7};
    assign wire1201 = {4'd9, 4'd7};
    assign wire1202 = {4'd9, 4'd7};
    assign wire1203 = {4'd9, 4'd7};
    assign wire1204 = {4'd10, 4'd8};
    assign wire1205 = {4'd9, 4'd7};
    assign wire1206 = {4'd9, 4'd7};
    assign wire1207 = {4'd9, 4'd7};
    assign wire1208 = {4'd5, 4'd3};
    assign wire1209 = {4'd5, 4'd3};
    assign wire1210 = {4'd5, 4'd3};
    assign wire1211 = {4'd5, 4'd3};
    assign wire1212 = {4'd5, 4'd3};
    assign wire1213 = {4'd5, 4'd3};
    assign wire1214 = {4'd5, 4'd3};
    assign wire1215 = {4'd5, 4'd3};
    assign wire1216 = {4'd7, 4'd3};
    assign wire1217 = {4'd7, 4'd3};
    assign wire1218 = {4'd7, 4'd3};
    assign wire1219 = {4'd7, 4'd3};
    assign wire1220 = {4'd8, 4'd4};
    assign wire1221 = {4'd11, 4'd7};
    assign wire1222 = {4'd7, 4'd3};
    assign wire1223 = {4'd7, 4'd3};
    assign wire1224 = {4'd8, 4'd4};
    assign wire1225 = {4'd8, 4'd4};
    assign wire1226 = {4'd8, 4'd4};
    assign wire1227 = {4'd8, 4'd4};
    assign wire1228 = {4'd9, 4'd5};
    assign wire1229 = {4'd8, 4'd4};
    assign wire1230 = {4'd8, 4'd4};
    assign wire1231 = {4'd8, 4'd4};
    assign wire1232 = {4'd11, 4'd7};
    assign wire1233 = {4'd11, 4'd7};
    assign wire1234 = {4'd11, 4'd7};
    assign wire1235 = {4'd11, 4'd7};
    assign wire1236 = {4'd12, 4'd8};
    assign wire1237 = {4'd11, 4'd7};
    assign wire1238 = {4'd11, 4'd7};
    assign wire1239 = {4'd11, 4'd7};
    assign wire1240 = {4'd7, 4'd3};
    assign wire1241 = {4'd7, 4'd3};
    assign wire1242 = {4'd7, 4'd3};
    assign wire1243 = {4'd7, 4'd3};
    assign wire1244 = {4'd7, 4'd3};
    assign wire1245 = {4'd7, 4'd3};
    assign wire1246 = {4'd7, 4'd3};
    assign wire1247 = {4'd7, 4'd3};
    assign wire1248 = {4'd9, 4'd3};
    assign wire1249 = {4'd9, 4'd3};
    assign wire1250 = {4'd9, 4'd3};
    assign wire1251 = {4'd9, 4'd3};
    assign wire1252 = {4'd10, 4'd4};
    assign wire1253 = {4'd13, 4'd7};
    assign wire1254 = {4'd9, 4'd3};
    assign wire1255 = {4'd9, 4'd3};
    assign wire1256 = {4'd10, 4'd4};
    assign wire1257 = {4'd10, 4'd4};
    assign wire1258 = {4'd10, 4'd4};
    assign wire1259 = {4'd10, 4'd4};
    assign wire1260 = {4'd11, 4'd5};
    assign wire1261 = {4'd10, 4'd4};
    assign wire1262 = {4'd10, 4'd4};
    assign wire1263 = {4'd10, 4'd4};
    assign wire1264 = {4'd13, 4'd7};
    assign wire1265 = {4'd13, 4'd7};
    assign wire1266 = {4'd13, 4'd7};
    assign wire1267 = {4'd13, 4'd7};
    assign wire1268 = {4'd14, 4'd8};
    assign wire1269 = {4'd13, 4'd7};
    assign wire1270 = {4'd13, 4'd7};
    assign wire1271 = {4'd13, 4'd7};
    assign wire1272 = {4'd9, 4'd3};
    assign wire1273 = {4'd9, 4'd3};
    assign wire1274 = {4'd9, 4'd3};
    assign wire1275 = {4'd9, 4'd3};
    assign wire1276 = {4'd9, 4'd3};
    assign wire1277 = {4'd9, 4'd3};
    assign wire1278 = {4'd9, 4'd3};
    assign wire1279 = {4'd9, 4'd3};
    assign wire1280 = {4'd4, 4'd3};
    assign wire1281 = {4'd4, 4'd3};
    assign wire1282 = {4'd4, 4'd3};
    assign wire1283 = {4'd4, 4'd3};
    assign wire1284 = {4'd4, 4'd3};
    assign wire1285 = {4'd4, 4'd3};
    assign wire1286 = {4'd4, 4'd3};
    assign wire1287 = {4'd4, 4'd3};
    assign wire1288 = {4'd4, 4'd3};
    assign wire1289 = {4'd4, 4'd3};
    assign wire1290 = {4'd4, 4'd3};
    assign wire1291 = {4'd4, 4'd3};
    assign wire1292 = {4'd4, 4'd3};
    assign wire1293 = {4'd4, 4'd3};
    assign wire1294 = {4'd4, 4'd3};
    assign wire1295 = {4'd4, 4'd3};
    assign wire1296 = {4'd4, 4'd3};
    assign wire1297 = {4'd4, 4'd3};
    assign wire1298 = {4'd4, 4'd3};
    assign wire1299 = {4'd4, 4'd3};
    assign wire1300 = {4'd4, 4'd3};
    assign wire1301 = {4'd4, 4'd3};
    assign wire1302 = {4'd4, 4'd3};
    assign wire1303 = {4'd4, 4'd3};
    assign wire1304 = {4'd4, 4'd3};
    assign wire1305 = {4'd4, 4'd3};
    assign wire1306 = {4'd4, 4'd3};
    assign wire1307 = {4'd4, 4'd3};
    assign wire1308 = {4'd4, 4'd3};
    assign wire1309 = {4'd4, 4'd3};
    assign wire1310 = {4'd4, 4'd3};
    assign wire1311 = {4'd4, 4'd3};
    assign wire1312 = {4'd5, 4'd3};
    assign wire1313 = {4'd5, 4'd3};
    assign wire1314 = {4'd5, 4'd3};
    assign wire1315 = {4'd5, 4'd3};
    assign wire1316 = {4'd5, 4'd3};
    assign wire1317 = {4'd5, 4'd3};
    assign wire1318 = {4'd5, 4'd3};
    assign wire1319 = {4'd5, 4'd3};
    assign wire1320 = {4'd5, 4'd3};
    assign wire1321 = {4'd5, 4'd3};
    assign wire1322 = {4'd5, 4'd3};
    assign wire1323 = {4'd5, 4'd3};
    assign wire1324 = {4'd5, 4'd3};
    assign wire1325 = {4'd5, 4'd3};
    assign wire1326 = {4'd5, 4'd3};
    assign wire1327 = {4'd5, 4'd3};
    assign wire1328 = {4'd5, 4'd3};
    assign wire1329 = {4'd5, 4'd3};
    assign wire1330 = {4'd5, 4'd3};
    assign wire1331 = {4'd5, 4'd3};
    assign wire1332 = {4'd5, 4'd3};
    assign wire1333 = {4'd5, 4'd3};
    assign wire1334 = {4'd5, 4'd3};
    assign wire1335 = {4'd5, 4'd3};
    assign wire1336 = {4'd5, 4'd3};
    assign wire1337 = {4'd5, 4'd3};
    assign wire1338 = {4'd5, 4'd3};
    assign wire1339 = {4'd5, 4'd3};
    assign wire1340 = {4'd5, 4'd3};
    assign wire1341 = {4'd5, 4'd3};
    assign wire1342 = {4'd5, 4'd3};
    assign wire1343 = {4'd5, 4'd3};
    assign wire1344 = {4'd7, 4'd3};
    assign wire1345 = {4'd7, 4'd3};
    assign wire1346 = {4'd7, 4'd3};
    assign wire1347 = {4'd7, 4'd3};
    assign wire1348 = {4'd7, 4'd3};
    assign wire1349 = {4'd7, 4'd3};
    assign wire1350 = {4'd7, 4'd3};
    assign wire1351 = {4'd7, 4'd3};
    assign wire1352 = {4'd7, 4'd3};
    assign wire1353 = {4'd7, 4'd3};
    assign wire1354 = {4'd7, 4'd3};
    assign wire1355 = {4'd7, 4'd3};
    assign wire1356 = {4'd7, 4'd3};
    assign wire1357 = {4'd7, 4'd3};
    assign wire1358 = {4'd7, 4'd3};
    assign wire1359 = {4'd7, 4'd3};
    assign wire1360 = {4'd7, 4'd3};
    assign wire1361 = {4'd7, 4'd3};
    assign wire1362 = {4'd7, 4'd3};
    assign wire1363 = {4'd7, 4'd3};
    assign wire1364 = {4'd7, 4'd3};
    assign wire1365 = {4'd7, 4'd3};
    assign wire1366 = {4'd7, 4'd3};
    assign wire1367 = {4'd7, 4'd3};
    assign wire1368 = {4'd7, 4'd3};
    assign wire1369 = {4'd7, 4'd3};
    assign wire1370 = {4'd7, 4'd3};
    assign wire1371 = {4'd7, 4'd3};
    assign wire1372 = {4'd7, 4'd3};
    assign wire1373 = {4'd7, 4'd3};
    assign wire1374 = {4'd7, 4'd3};
    assign wire1375 = {4'd7, 4'd3};
    assign wire1376 = {4'd9, 4'd3};
    assign wire1377 = {4'd9, 4'd3};
    assign wire1378 = {4'd9, 4'd3};
    assign wire1379 = {4'd9, 4'd3};
    assign wire1380 = {4'd9, 4'd3};
    assign wire1381 = {4'd9, 4'd3};
    assign wire1382 = {4'd9, 4'd3};
    assign wire1383 = {4'd9, 4'd3};
    assign wire1384 = {4'd9, 4'd3};
    assign wire1385 = {4'd9, 4'd3};
    assign wire1386 = {4'd9, 4'd3};
    assign wire1387 = {4'd9, 4'd3};
    assign wire1388 = {4'd9, 4'd3};
    assign wire1389 = {4'd9, 4'd3};
    assign wire1390 = {4'd9, 4'd3};
    assign wire1391 = {4'd9, 4'd3};
    assign wire1392 = {4'd9, 4'd3};
    assign wire1393 = {4'd9, 4'd3};
    assign wire1394 = {4'd9, 4'd3};
    assign wire1395 = {4'd9, 4'd3};
    assign wire1396 = {4'd9, 4'd3};
    assign wire1397 = {4'd9, 4'd3};
    assign wire1398 = {4'd9, 4'd3};
    assign wire1399 = {4'd9, 4'd3};
    assign wire1400 = {4'd9, 4'd3};
    assign wire1401 = {4'd9, 4'd3};
    assign wire1402 = {4'd9, 4'd3};
    assign wire1403 = {4'd9, 4'd3};
    assign wire1404 = {4'd9, 4'd3};
    assign wire1405 = {4'd9, 4'd3};
    assign wire1406 = {4'd9, 4'd3};
    assign wire1407 = {4'd9, 4'd3};
    assign wire1408 = {4'd5, 4'd4};
    assign wire1409 = {4'd5, 4'd4};
    assign wire1410 = {4'd5, 4'd4};
    assign wire1411 = {4'd5, 4'd4};
    assign wire1412 = {4'd6, 4'd5};
    assign wire1413 = {4'd9, 4'd8};
    assign wire1414 = {4'd5, 4'd4};
    assign wire1415 = {4'd5, 4'd4};
    assign wire1416 = {4'd6, 4'd5};
    assign wire1417 = {4'd6, 4'd5};
    assign wire1418 = {4'd6, 4'd5};
    assign wire1419 = {4'd6, 4'd5};
    assign wire1420 = {4'd7, 4'd6};
    assign wire1421 = {4'd6, 4'd5};
    assign wire1422 = {4'd6, 4'd5};
    assign wire1423 = {4'd6, 4'd5};
    assign wire1424 = {4'd9, 4'd8};
    assign wire1425 = {4'd9, 4'd8};
    assign wire1426 = {4'd9, 4'd8};
    assign wire1427 = {4'd9, 4'd8};
    assign wire1428 = {4'd10, 4'd9};
    assign wire1429 = {4'd9, 4'd8};
    assign wire1430 = {4'd9, 4'd8};
    assign wire1431 = {4'd9, 4'd8};
    assign wire1432 = {4'd5, 4'd4};
    assign wire1433 = {4'd5, 4'd4};
    assign wire1434 = {4'd5, 4'd4};
    assign wire1435 = {4'd5, 4'd4};
    assign wire1436 = {4'd5, 4'd4};
    assign wire1437 = {4'd5, 4'd4};
    assign wire1438 = {4'd5, 4'd4};
    assign wire1439 = {4'd5, 4'd4};
    assign wire1440 = {4'd6, 4'd4};
    assign wire1441 = {4'd6, 4'd4};
    assign wire1442 = {4'd6, 4'd4};
    assign wire1443 = {4'd6, 4'd4};
    assign wire1444 = {4'd7, 4'd5};
    assign wire1445 = {4'd10, 4'd8};
    assign wire1446 = {4'd6, 4'd4};
    assign wire1447 = {4'd6, 4'd4};
    assign wire1448 = {4'd7, 4'd5};
    assign wire1449 = {4'd7, 4'd5};
    assign wire1450 = {4'd7, 4'd5};
    assign wire1451 = {4'd7, 4'd5};
    assign wire1452 = {4'd8, 4'd6};
    assign wire1453 = {4'd7, 4'd5};
    assign wire1454 = {4'd7, 4'd5};
    assign wire1455 = {4'd7, 4'd5};
    assign wire1456 = {4'd10, 4'd8};
    assign wire1457 = {4'd10, 4'd8};
    assign wire1458 = {4'd10, 4'd8};
    assign wire1459 = {4'd10, 4'd8};
    assign wire1460 = {4'd11, 4'd9};
    assign wire1461 = {4'd10, 4'd8};
    assign wire1462 = {4'd10, 4'd8};
    assign wire1463 = {4'd10, 4'd8};
    assign wire1464 = {4'd6, 4'd4};
    assign wire1465 = {4'd6, 4'd4};
    assign wire1466 = {4'd6, 4'd4};
    assign wire1467 = {4'd6, 4'd4};
    assign wire1468 = {4'd6, 4'd4};
    assign wire1469 = {4'd6, 4'd4};
    assign wire1470 = {4'd6, 4'd4};
    assign wire1471 = {4'd6, 4'd4};
    assign wire1472 = {4'd8, 4'd4};
    assign wire1473 = {4'd8, 4'd4};
    assign wire1474 = {4'd8, 4'd4};
    assign wire1475 = {4'd8, 4'd4};
    assign wire1476 = {4'd9, 4'd5};
    assign wire1477 = {4'd12, 4'd8};
    assign wire1478 = {4'd8, 4'd4};
    assign wire1479 = {4'd8, 4'd4};
    assign wire1480 = {4'd9, 4'd5};
    assign wire1481 = {4'd9, 4'd5};
    assign wire1482 = {4'd9, 4'd5};
    assign wire1483 = {4'd9, 4'd5};
    assign wire1484 = {4'd10, 4'd6};
    assign wire1485 = {4'd9, 4'd5};
    assign wire1486 = {4'd9, 4'd5};
    assign wire1487 = {4'd9, 4'd5};
    assign wire1488 = {4'd12, 4'd8};
    assign wire1489 = {4'd12, 4'd8};
    assign wire1490 = {4'd12, 4'd8};
    assign wire1491 = {4'd12, 4'd8};
    assign wire1492 = {4'd13, 4'd9};
    assign wire1493 = {4'd12, 4'd8};
    assign wire1494 = {4'd12, 4'd8};
    assign wire1495 = {4'd12, 4'd8};
    assign wire1496 = {4'd8, 4'd4};
    assign wire1497 = {4'd8, 4'd4};
    assign wire1498 = {4'd8, 4'd4};
    assign wire1499 = {4'd8, 4'd4};
    assign wire1500 = {4'd8, 4'd4};
    assign wire1501 = {4'd8, 4'd4};
    assign wire1502 = {4'd8, 4'd4};
    assign wire1503 = {4'd8, 4'd4};
    assign wire1504 = {4'd10, 4'd4};
    assign wire1505 = {4'd10, 4'd4};
    assign wire1506 = {4'd10, 4'd4};
    assign wire1507 = {4'd10, 4'd4};
    assign wire1508 = {4'd11, 4'd5};
    assign wire1509 = {4'd14, 4'd8};
    assign wire1510 = {4'd10, 4'd4};
    assign wire1511 = {4'd10, 4'd4};
    assign wire1512 = {4'd11, 4'd5};
    assign wire1513 = {4'd11, 4'd5};
    assign wire1514 = {4'd11, 4'd5};
    assign wire1515 = {4'd11, 4'd5};
    assign wire1516 = {4'd12, 4'd6};
    assign wire1517 = {4'd11, 4'd5};
    assign wire1518 = {4'd11, 4'd5};
    assign wire1519 = {4'd11, 4'd5};
    assign wire1520 = {4'd14, 4'd8};
    assign wire1521 = {4'd14, 4'd8};
    assign wire1522 = {4'd14, 4'd8};
    assign wire1523 = {4'd14, 4'd8};
    assign wire1524 = {4'd15, 4'd9};
    assign wire1525 = {4'd14, 4'd8};
    assign wire1526 = {4'd14, 4'd8};
    assign wire1527 = {4'd14, 4'd8};
    assign wire1528 = {4'd10, 4'd4};
    assign wire1529 = {4'd10, 4'd4};
    assign wire1530 = {4'd10, 4'd4};
    assign wire1531 = {4'd10, 4'd4};
    assign wire1532 = {4'd10, 4'd4};
    assign wire1533 = {4'd10, 4'd4};
    assign wire1534 = {4'd10, 4'd4};
    assign wire1535 = {4'd10, 4'd4};
    assign wire1536 = {4'd4, 4'd3};
    assign wire1537 = {4'd4, 4'd3};
    assign wire1538 = {4'd4, 4'd3};
    assign wire1539 = {4'd4, 4'd3};
    assign wire1540 = {4'd4, 4'd3};
    assign wire1541 = {4'd4, 4'd3};
    assign wire1542 = {4'd4, 4'd3};
    assign wire1543 = {4'd4, 4'd3};
    assign wire1544 = {4'd4, 4'd3};
    assign wire1545 = {4'd4, 4'd3};
    assign wire1546 = {4'd4, 4'd3};
    assign wire1547 = {4'd4, 4'd3};
    assign wire1548 = {4'd4, 4'd3};
    assign wire1549 = {4'd4, 4'd3};
    assign wire1550 = {4'd4, 4'd3};
    assign wire1551 = {4'd4, 4'd3};
    assign wire1552 = {4'd4, 4'd3};
    assign wire1553 = {4'd4, 4'd3};
    assign wire1554 = {4'd4, 4'd3};
    assign wire1555 = {4'd4, 4'd3};
    assign wire1556 = {4'd4, 4'd3};
    assign wire1557 = {4'd4, 4'd3};
    assign wire1558 = {4'd4, 4'd3};
    assign wire1559 = {4'd4, 4'd3};
    assign wire1560 = {4'd4, 4'd3};
    assign wire1561 = {4'd4, 4'd3};
    assign wire1562 = {4'd4, 4'd3};
    assign wire1563 = {4'd4, 4'd3};
    assign wire1564 = {4'd4, 4'd3};
    assign wire1565 = {4'd4, 4'd3};
    assign wire1566 = {4'd4, 4'd3};
    assign wire1567 = {4'd4, 4'd3};
    assign wire1568 = {4'd5, 4'd3};
    assign wire1569 = {4'd5, 4'd3};
    assign wire1570 = {4'd5, 4'd3};
    assign wire1571 = {4'd5, 4'd3};
    assign wire1572 = {4'd5, 4'd3};
    assign wire1573 = {4'd5, 4'd3};
    assign wire1574 = {4'd5, 4'd3};
    assign wire1575 = {4'd5, 4'd3};
    assign wire1576 = {4'd5, 4'd3};
    assign wire1577 = {4'd5, 4'd3};
    assign wire1578 = {4'd5, 4'd3};
    assign wire1579 = {4'd5, 4'd3};
    assign wire1580 = {4'd5, 4'd3};
    assign wire1581 = {4'd5, 4'd3};
    assign wire1582 = {4'd5, 4'd3};
    assign wire1583 = {4'd5, 4'd3};
    assign wire1584 = {4'd5, 4'd3};
    assign wire1585 = {4'd5, 4'd3};
    assign wire1586 = {4'd5, 4'd3};
    assign wire1587 = {4'd5, 4'd3};
    assign wire1588 = {4'd5, 4'd3};
    assign wire1589 = {4'd5, 4'd3};
    assign wire1590 = {4'd5, 4'd3};
    assign wire1591 = {4'd5, 4'd3};
    assign wire1592 = {4'd5, 4'd3};
    assign wire1593 = {4'd5, 4'd3};
    assign wire1594 = {4'd5, 4'd3};
    assign wire1595 = {4'd5, 4'd3};
    assign wire1596 = {4'd5, 4'd3};
    assign wire1597 = {4'd5, 4'd3};
    assign wire1598 = {4'd5, 4'd3};
    assign wire1599 = {4'd5, 4'd3};
    assign wire1600 = {4'd7, 4'd3};
    assign wire1601 = {4'd7, 4'd3};
    assign wire1602 = {4'd7, 4'd3};
    assign wire1603 = {4'd7, 4'd3};
    assign wire1604 = {4'd7, 4'd3};
    assign wire1605 = {4'd7, 4'd3};
    assign wire1606 = {4'd7, 4'd3};
    assign wire1607 = {4'd7, 4'd3};
    assign wire1608 = {4'd7, 4'd3};
    assign wire1609 = {4'd7, 4'd3};
    assign wire1610 = {4'd7, 4'd3};
    assign wire1611 = {4'd7, 4'd3};
    assign wire1612 = {4'd7, 4'd3};
    assign wire1613 = {4'd7, 4'd3};
    assign wire1614 = {4'd7, 4'd3};
    assign wire1615 = {4'd7, 4'd3};
    assign wire1616 = {4'd7, 4'd3};
    assign wire1617 = {4'd7, 4'd3};
    assign wire1618 = {4'd7, 4'd3};
    assign wire1619 = {4'd7, 4'd3};
    assign wire1620 = {4'd7, 4'd3};
    assign wire1621 = {4'd7, 4'd3};
    assign wire1622 = {4'd7, 4'd3};
    assign wire1623 = {4'd7, 4'd3};
    assign wire1624 = {4'd7, 4'd3};
    assign wire1625 = {4'd7, 4'd3};
    assign wire1626 = {4'd7, 4'd3};
    assign wire1627 = {4'd7, 4'd3};
    assign wire1628 = {4'd7, 4'd3};
    assign wire1629 = {4'd7, 4'd3};
    assign wire1630 = {4'd7, 4'd3};
    assign wire1631 = {4'd7, 4'd3};
    assign wire1632 = {4'd9, 4'd3};
    assign wire1633 = {4'd9, 4'd3};
    assign wire1634 = {4'd9, 4'd3};
    assign wire1635 = {4'd9, 4'd3};
    assign wire1636 = {4'd9, 4'd3};
    assign wire1637 = {4'd9, 4'd3};
    assign wire1638 = {4'd9, 4'd3};
    assign wire1639 = {4'd9, 4'd3};
    assign wire1640 = {4'd9, 4'd3};
    assign wire1641 = {4'd9, 4'd3};
    assign wire1642 = {4'd9, 4'd3};
    assign wire1643 = {4'd9, 4'd3};
    assign wire1644 = {4'd9, 4'd3};
    assign wire1645 = {4'd9, 4'd3};
    assign wire1646 = {4'd9, 4'd3};
    assign wire1647 = {4'd9, 4'd3};
    assign wire1648 = {4'd9, 4'd3};
    assign wire1649 = {4'd9, 4'd3};
    assign wire1650 = {4'd9, 4'd3};
    assign wire1651 = {4'd9, 4'd3};
    assign wire1652 = {4'd9, 4'd3};
    assign wire1653 = {4'd9, 4'd3};
    assign wire1654 = {4'd9, 4'd3};
    assign wire1655 = {4'd9, 4'd3};
    assign wire1656 = {4'd9, 4'd3};
    assign wire1657 = {4'd9, 4'd3};
    assign wire1658 = {4'd9, 4'd3};
    assign wire1659 = {4'd9, 4'd3};
    assign wire1660 = {4'd9, 4'd3};
    assign wire1661 = {4'd9, 4'd3};
    assign wire1662 = {4'd9, 4'd3};
    assign wire1663 = {4'd9, 4'd3};
    assign wire1664 = {4'd5, 4'd4};
    assign wire1665 = {4'd5, 4'd4};
    assign wire1666 = {4'd5, 4'd4};
    assign wire1667 = {4'd5, 4'd4};
    assign wire1668 = {4'd5, 4'd4};
    assign wire1669 = {4'd7, 4'd6};
    assign wire1670 = {4'd5, 4'd4};
    assign wire1671 = {4'd5, 4'd4};
    assign wire1672 = {4'd6, 4'd5};
    assign wire1673 = {4'd6, 4'd5};
    assign wire1674 = {4'd6, 4'd5};
    assign wire1675 = {4'd6, 4'd5};
    assign wire1676 = {4'd6, 4'd5};
    assign wire1677 = {4'd6, 4'd5};
    assign wire1678 = {4'd6, 4'd5};
    assign wire1679 = {4'd6, 4'd5};
    assign wire1680 = {4'd7, 4'd6};
    assign wire1681 = {4'd7, 4'd6};
    assign wire1682 = {4'd7, 4'd6};
    assign wire1683 = {4'd7, 4'd6};
    assign wire1684 = {4'd7, 4'd6};
    assign wire1685 = {4'd7, 4'd6};
    assign wire1686 = {4'd7, 4'd6};
    assign wire1687 = {4'd7, 4'd6};
    assign wire1688 = {4'd5, 4'd4};
    assign wire1689 = {4'd5, 4'd4};
    assign wire1690 = {4'd5, 4'd4};
    assign wire1691 = {4'd5, 4'd4};
    assign wire1692 = {4'd5, 4'd4};
    assign wire1693 = {4'd5, 4'd4};
    assign wire1694 = {4'd5, 4'd4};
    assign wire1695 = {4'd5, 4'd4};
    assign wire1696 = {4'd6, 4'd4};
    assign wire1697 = {4'd6, 4'd4};
    assign wire1698 = {4'd6, 4'd4};
    assign wire1699 = {4'd6, 4'd4};
    assign wire1700 = {4'd6, 4'd4};
    assign wire1701 = {4'd8, 4'd6};
    assign wire1702 = {4'd6, 4'd4};
    assign wire1703 = {4'd6, 4'd4};
    assign wire1704 = {4'd7, 4'd5};
    assign wire1705 = {4'd7, 4'd5};
    assign wire1706 = {4'd7, 4'd5};
    assign wire1707 = {4'd7, 4'd5};
    assign wire1708 = {4'd7, 4'd5};
    assign wire1709 = {4'd7, 4'd5};
    assign wire1710 = {4'd7, 4'd5};
    assign wire1711 = {4'd7, 4'd5};
    assign wire1712 = {4'd8, 4'd6};
    assign wire1713 = {4'd8, 4'd6};
    assign wire1714 = {4'd8, 4'd6};
    assign wire1715 = {4'd8, 4'd6};
    assign wire1716 = {4'd8, 4'd6};
    assign wire1717 = {4'd8, 4'd6};
    assign wire1718 = {4'd8, 4'd6};
    assign wire1719 = {4'd8, 4'd6};
    assign wire1720 = {4'd6, 4'd4};
    assign wire1721 = {4'd6, 4'd4};
    assign wire1722 = {4'd6, 4'd4};
    assign wire1723 = {4'd6, 4'd4};
    assign wire1724 = {4'd6, 4'd4};
    assign wire1725 = {4'd6, 4'd4};
    assign wire1726 = {4'd6, 4'd4};
    assign wire1727 = {4'd6, 4'd4};
    assign wire1728 = {4'd8, 4'd4};
    assign wire1729 = {4'd8, 4'd4};
    assign wire1730 = {4'd8, 4'd4};
    assign wire1731 = {4'd8, 4'd4};
    assign wire1732 = {4'd8, 4'd4};
    assign wire1733 = {4'd10, 4'd6};
    assign wire1734 = {4'd8, 4'd4};
    assign wire1735 = {4'd8, 4'd4};
    assign wire1736 = {4'd9, 4'd5};
    assign wire1737 = {4'd9, 4'd5};
    assign wire1738 = {4'd9, 4'd5};
    assign wire1739 = {4'd9, 4'd5};
    assign wire1740 = {4'd9, 4'd5};
    assign wire1741 = {4'd9, 4'd5};
    assign wire1742 = {4'd9, 4'd5};
    assign wire1743 = {4'd9, 4'd5};
    assign wire1744 = {4'd10, 4'd6};
    assign wire1745 = {4'd10, 4'd6};
    assign wire1746 = {4'd10, 4'd6};
    assign wire1747 = {4'd10, 4'd6};
    assign wire1748 = {4'd10, 4'd6};
    assign wire1749 = {4'd10, 4'd6};
    assign wire1750 = {4'd10, 4'd6};
    assign wire1751 = {4'd10, 4'd6};
    assign wire1752 = {4'd8, 4'd4};
    assign wire1753 = {4'd8, 4'd4};
    assign wire1754 = {4'd8, 4'd4};
    assign wire1755 = {4'd8, 4'd4};
    assign wire1756 = {4'd8, 4'd4};
    assign wire1757 = {4'd8, 4'd4};
    assign wire1758 = {4'd8, 4'd4};
    assign wire1759 = {4'd8, 4'd4};
    assign wire1760 = {4'd10, 4'd4};
    assign wire1761 = {4'd10, 4'd4};
    assign wire1762 = {4'd10, 4'd4};
    assign wire1763 = {4'd10, 4'd4};
    assign wire1764 = {4'd10, 4'd4};
    assign wire1765 = {4'd12, 4'd6};
    assign wire1766 = {4'd10, 4'd4};
    assign wire1767 = {4'd10, 4'd4};
    assign wire1768 = {4'd11, 4'd5};
    assign wire1769 = {4'd11, 4'd5};
    assign wire1770 = {4'd11, 4'd5};
    assign wire1771 = {4'd11, 4'd5};
    assign wire1772 = {4'd11, 4'd5};
    assign wire1773 = {4'd11, 4'd5};
    assign wire1774 = {4'd11, 4'd5};
    assign wire1775 = {4'd11, 4'd5};
    assign wire1776 = {4'd12, 4'd6};
    assign wire1777 = {4'd12, 4'd6};
    assign wire1778 = {4'd12, 4'd6};
    assign wire1779 = {4'd12, 4'd6};
    assign wire1780 = {4'd12, 4'd6};
    assign wire1781 = {4'd12, 4'd6};
    assign wire1782 = {4'd12, 4'd6};
    assign wire1783 = {4'd12, 4'd6};
    assign wire1784 = {4'd10, 4'd4};
    assign wire1785 = {4'd10, 4'd4};
    assign wire1786 = {4'd10, 4'd4};
    assign wire1787 = {4'd10, 4'd4};
    assign wire1788 = {4'd10, 4'd4};
    assign wire1789 = {4'd10, 4'd4};
    assign wire1790 = {4'd10, 4'd4};
    assign wire1791 = {4'd10, 4'd4};
    assign wire1792 = {4'd5, 4'd4};
    assign wire1793 = {4'd5, 4'd4};
    assign wire1794 = {4'd5, 4'd4};
    assign wire1795 = {4'd5, 4'd4};
    assign wire1796 = {4'd5, 4'd4};
    assign wire1797 = {4'd5, 4'd4};
    assign wire1798 = {4'd5, 4'd4};
    assign wire1799 = {4'd5, 4'd4};
    assign wire1800 = {4'd5, 4'd4};
    assign wire1801 = {4'd5, 4'd4};
    assign wire1802 = {4'd5, 4'd4};
    assign wire1803 = {4'd5, 4'd4};
    assign wire1804 = {4'd5, 4'd4};
    assign wire1805 = {4'd5, 4'd4};
    assign wire1806 = {4'd5, 4'd4};
    assign wire1807 = {4'd5, 4'd4};
    assign wire1808 = {4'd5, 4'd4};
    assign wire1809 = {4'd5, 4'd4};
    assign wire1810 = {4'd5, 4'd4};
    assign wire1811 = {4'd5, 4'd4};
    assign wire1812 = {4'd5, 4'd4};
    assign wire1813 = {4'd5, 4'd4};
    assign wire1814 = {4'd5, 4'd4};
    assign wire1815 = {4'd5, 4'd4};
    assign wire1816 = {4'd5, 4'd4};
    assign wire1817 = {4'd5, 4'd4};
    assign wire1818 = {4'd5, 4'd4};
    assign wire1819 = {4'd5, 4'd4};
    assign wire1820 = {4'd5, 4'd4};
    assign wire1821 = {4'd5, 4'd4};
    assign wire1822 = {4'd5, 4'd4};
    assign wire1823 = {4'd5, 4'd4};
    assign wire1824 = {4'd6, 4'd4};
    assign wire1825 = {4'd6, 4'd4};
    assign wire1826 = {4'd6, 4'd4};
    assign wire1827 = {4'd6, 4'd4};
    assign wire1828 = {4'd6, 4'd4};
    assign wire1829 = {4'd6, 4'd4};
    assign wire1830 = {4'd6, 4'd4};
    assign wire1831 = {4'd6, 4'd4};
    assign wire1832 = {4'd6, 4'd4};
    assign wire1833 = {4'd6, 4'd4};
    assign wire1834 = {4'd6, 4'd4};
    assign wire1835 = {4'd6, 4'd4};
    assign wire1836 = {4'd6, 4'd4};
    assign wire1837 = {4'd6, 4'd4};
    assign wire1838 = {4'd6, 4'd4};
    assign wire1839 = {4'd6, 4'd4};
    assign wire1840 = {4'd6, 4'd4};
    assign wire1841 = {4'd6, 4'd4};
    assign wire1842 = {4'd6, 4'd4};
    assign wire1843 = {4'd6, 4'd4};
    assign wire1844 = {4'd6, 4'd4};
    assign wire1845 = {4'd6, 4'd4};
    assign wire1846 = {4'd6, 4'd4};
    assign wire1847 = {4'd6, 4'd4};
    assign wire1848 = {4'd6, 4'd4};
    assign wire1849 = {4'd6, 4'd4};
    assign wire1850 = {4'd6, 4'd4};
    assign wire1851 = {4'd6, 4'd4};
    assign wire1852 = {4'd6, 4'd4};
    assign wire1853 = {4'd6, 4'd4};
    assign wire1854 = {4'd6, 4'd4};
    assign wire1855 = {4'd6, 4'd4};
    assign wire1856 = {4'd8, 4'd4};
    assign wire1857 = {4'd8, 4'd4};
    assign wire1858 = {4'd8, 4'd4};
    assign wire1859 = {4'd8, 4'd4};
    assign wire1860 = {4'd8, 4'd4};
    assign wire1861 = {4'd8, 4'd4};
    assign wire1862 = {4'd8, 4'd4};
    assign wire1863 = {4'd8, 4'd4};
    assign wire1864 = {4'd8, 4'd4};
    assign wire1865 = {4'd8, 4'd4};
    assign wire1866 = {4'd8, 4'd4};
    assign wire1867 = {4'd8, 4'd4};
    assign wire1868 = {4'd8, 4'd4};
    assign wire1869 = {4'd8, 4'd4};
    assign wire1870 = {4'd8, 4'd4};
    assign wire1871 = {4'd8, 4'd4};
    assign wire1872 = {4'd8, 4'd4};
    assign wire1873 = {4'd8, 4'd4};
    assign wire1874 = {4'd8, 4'd4};
    assign wire1875 = {4'd8, 4'd4};
    assign wire1876 = {4'd8, 4'd4};
    assign wire1877 = {4'd8, 4'd4};
    assign wire1878 = {4'd8, 4'd4};
    assign wire1879 = {4'd8, 4'd4};
    assign wire1880 = {4'd8, 4'd4};
    assign wire1881 = {4'd8, 4'd4};
    assign wire1882 = {4'd8, 4'd4};
    assign wire1883 = {4'd8, 4'd4};
    assign wire1884 = {4'd8, 4'd4};
    assign wire1885 = {4'd8, 4'd4};
    assign wire1886 = {4'd8, 4'd4};
    assign wire1887 = {4'd8, 4'd4};
    assign wire1888 = {4'd10, 4'd4};
    assign wire1889 = {4'd10, 4'd4};
    assign wire1890 = {4'd10, 4'd4};
    assign wire1891 = {4'd10, 4'd4};
    assign wire1892 = {4'd10, 4'd4};
    assign wire1893 = {4'd10, 4'd4};
    assign wire1894 = {4'd10, 4'd4};
    assign wire1895 = {4'd10, 4'd4};
    assign wire1896 = {4'd10, 4'd4};
    assign wire1897 = {4'd10, 4'd4};
    assign wire1898 = {4'd10, 4'd4};
    assign wire1899 = {4'd10, 4'd4};
    assign wire1900 = {4'd10, 4'd4};
    assign wire1901 = {4'd10, 4'd4};
    assign wire1902 = {4'd10, 4'd4};
    assign wire1903 = {4'd10, 4'd4};
    assign wire1904 = {4'd10, 4'd4};
    assign wire1905 = {4'd10, 4'd4};
    assign wire1906 = {4'd10, 4'd4};
    assign wire1907 = {4'd10, 4'd4};
    assign wire1908 = {4'd10, 4'd4};
    assign wire1909 = {4'd10, 4'd4};
    assign wire1910 = {4'd10, 4'd4};
    assign wire1911 = {4'd10, 4'd4};
    assign wire1912 = {4'd10, 4'd4};
    assign wire1913 = {4'd10, 4'd4};
    assign wire1914 = {4'd10, 4'd4};
    assign wire1915 = {4'd10, 4'd4};
    assign wire1916 = {4'd10, 4'd4};
    assign wire1917 = {4'd10, 4'd4};
    assign wire1918 = {4'd10, 4'd4};
    assign wire1919 = {4'd10, 4'd4};
    assign wire1920 = {4'd6, 4'd5};
    assign wire1921 = {4'd6, 4'd5};
    assign wire1922 = {4'd6, 4'd5};
    assign wire1923 = {4'd6, 4'd5};
    assign wire1924 = {4'd6, 4'd5};
    assign wire1925 = {4'd8, 4'd7};
    assign wire1926 = {4'd6, 4'd5};
    assign wire1927 = {4'd6, 4'd5};
    assign wire1928 = {4'd7, 4'd6};
    assign wire1929 = {4'd7, 4'd6};
    assign wire1930 = {4'd7, 4'd6};
    assign wire1931 = {4'd7, 4'd6};
    assign wire1932 = {4'd7, 4'd6};
    assign wire1933 = {4'd7, 4'd6};
    assign wire1934 = {4'd7, 4'd6};
    assign wire1935 = {4'd7, 4'd6};
    assign wire1936 = {4'd8, 4'd7};
    assign wire1937 = {4'd8, 4'd7};
    assign wire1938 = {4'd8, 4'd7};
    assign wire1939 = {4'd8, 4'd7};
    assign wire1940 = {4'd8, 4'd7};
    assign wire1941 = {4'd8, 4'd7};
    assign wire1942 = {4'd8, 4'd7};
    assign wire1943 = {4'd8, 4'd7};
    assign wire1944 = {4'd6, 4'd5};
    assign wire1945 = {4'd6, 4'd5};
    assign wire1946 = {4'd6, 4'd5};
    assign wire1947 = {4'd6, 4'd5};
    assign wire1948 = {4'd6, 4'd5};
    assign wire1949 = {4'd6, 4'd5};
    assign wire1950 = {4'd6, 4'd5};
    assign wire1951 = {4'd6, 4'd5};
    assign wire1952 = {4'd7, 4'd5};
    assign wire1953 = {4'd7, 4'd5};
    assign wire1954 = {4'd7, 4'd5};
    assign wire1955 = {4'd7, 4'd5};
    assign wire1956 = {4'd7, 4'd5};
    assign wire1957 = {4'd9, 4'd7};
    assign wire1958 = {4'd7, 4'd5};
    assign wire1959 = {4'd7, 4'd5};
    assign wire1960 = {4'd8, 4'd6};
    assign wire1961 = {4'd8, 4'd6};
    assign wire1962 = {4'd8, 4'd6};
    assign wire1963 = {4'd8, 4'd6};
    assign wire1964 = {4'd8, 4'd6};
    assign wire1965 = {4'd8, 4'd6};
    assign wire1966 = {4'd8, 4'd6};
    assign wire1967 = {4'd8, 4'd6};
    assign wire1968 = {4'd9, 4'd7};
    assign wire1969 = {4'd9, 4'd7};
    assign wire1970 = {4'd9, 4'd7};
    assign wire1971 = {4'd9, 4'd7};
    assign wire1972 = {4'd9, 4'd7};
    assign wire1973 = {4'd9, 4'd7};
    assign wire1974 = {4'd9, 4'd7};
    assign wire1975 = {4'd9, 4'd7};
    assign wire1976 = {4'd7, 4'd5};
    assign wire1977 = {4'd7, 4'd5};
    assign wire1978 = {4'd7, 4'd5};
    assign wire1979 = {4'd7, 4'd5};
    assign wire1980 = {4'd7, 4'd5};
    assign wire1981 = {4'd7, 4'd5};
    assign wire1982 = {4'd7, 4'd5};
    assign wire1983 = {4'd7, 4'd5};
    assign wire1984 = {4'd9, 4'd5};
    assign wire1985 = {4'd9, 4'd5};
    assign wire1986 = {4'd9, 4'd5};
    assign wire1987 = {4'd9, 4'd5};
    assign wire1988 = {4'd9, 4'd5};
    assign wire1989 = {4'd11, 4'd7};
    assign wire1990 = {4'd9, 4'd5};
    assign wire1991 = {4'd9, 4'd5};
    assign wire1992 = {4'd10, 4'd6};
    assign wire1993 = {4'd10, 4'd6};
    assign wire1994 = {4'd10, 4'd6};
    assign wire1995 = {4'd10, 4'd6};
    assign wire1996 = {4'd10, 4'd6};
    assign wire1997 = {4'd10, 4'd6};
    assign wire1998 = {4'd10, 4'd6};
    assign wire1999 = {4'd10, 4'd6};
    assign wire2000 = {4'd11, 4'd7};
    assign wire2001 = {4'd11, 4'd7};
    assign wire2002 = {4'd11, 4'd7};
    assign wire2003 = {4'd11, 4'd7};
    assign wire2004 = {4'd11, 4'd7};
    assign wire2005 = {4'd11, 4'd7};
    assign wire2006 = {4'd11, 4'd7};
    assign wire2007 = {4'd11, 4'd7};
    assign wire2008 = {4'd9, 4'd5};
    assign wire2009 = {4'd9, 4'd5};
    assign wire2010 = {4'd9, 4'd5};
    assign wire2011 = {4'd9, 4'd5};
    assign wire2012 = {4'd9, 4'd5};
    assign wire2013 = {4'd9, 4'd5};
    assign wire2014 = {4'd9, 4'd5};
    assign wire2015 = {4'd9, 4'd5};
    assign wire2016 = {4'd11, 4'd5};
    assign wire2017 = {4'd11, 4'd5};
    assign wire2018 = {4'd11, 4'd5};
    assign wire2019 = {4'd11, 4'd5};
    assign wire2020 = {4'd11, 4'd5};
    assign wire2021 = {4'd13, 4'd7};
    assign wire2022 = {4'd11, 4'd5};
    assign wire2023 = {4'd11, 4'd5};
    assign wire2024 = {4'd12, 4'd6};
    assign wire2025 = {4'd12, 4'd6};
    assign wire2026 = {4'd12, 4'd6};
    assign wire2027 = {4'd12, 4'd6};
    assign wire2028 = {4'd12, 4'd6};
    assign wire2029 = {4'd12, 4'd6};
    assign wire2030 = {4'd12, 4'd6};
    assign wire2031 = {4'd12, 4'd6};
    assign wire2032 = {4'd13, 4'd7};
    assign wire2033 = {4'd13, 4'd7};
    assign wire2034 = {4'd13, 4'd7};
    assign wire2035 = {4'd13, 4'd7};
    assign wire2036 = {4'd13, 4'd7};
    assign wire2037 = {4'd13, 4'd7};
    assign wire2038 = {4'd13, 4'd7};
    assign wire2039 = {4'd13, 4'd7};
    assign wire2040 = {4'd11, 4'd5};
    assign wire2041 = {4'd11, 4'd5};
    assign wire2042 = {4'd11, 4'd5};
    assign wire2043 = {4'd11, 4'd5};
    assign wire2044 = {4'd11, 4'd5};
    assign wire2045 = {4'd11, 4'd5};
    assign wire2046 = {4'd11, 4'd5};
    assign wire2047 = {4'd11, 4'd5};
    assign wire2048 = {4'd3, 4'd2};
    assign wire2049 = {4'd3, 4'd2};
    assign wire2050 = {4'd3, 4'd2};
    assign wire2051 = {4'd3, 4'd2};
    assign wire2052 = {4'd3, 4'd2};
    assign wire2053 = {4'd3, 4'd2};
    assign wire2054 = {4'd3, 4'd2};
    assign wire2055 = {4'd3, 4'd2};
    assign wire2056 = {4'd3, 4'd2};
    assign wire2057 = {4'd3, 4'd2};
    assign wire2058 = {4'd3, 4'd2};
    assign wire2059 = {4'd3, 4'd2};
    assign wire2060 = {4'd3, 4'd2};
    assign wire2061 = {4'd3, 4'd2};
    assign wire2062 = {4'd3, 4'd2};
    assign wire2063 = {4'd3, 4'd2};
    assign wire2064 = {4'd3, 4'd2};
    assign wire2065 = {4'd3, 4'd2};
    assign wire2066 = {4'd3, 4'd2};
    assign wire2067 = {4'd3, 4'd2};
    assign wire2068 = {4'd3, 4'd2};
    assign wire2069 = {4'd3, 4'd2};
    assign wire2070 = {4'd3, 4'd2};
    assign wire2071 = {4'd3, 4'd2};
    assign wire2072 = {4'd3, 4'd2};
    assign wire2073 = {4'd3, 4'd2};
    assign wire2074 = {4'd3, 4'd2};
    assign wire2075 = {4'd3, 4'd2};
    assign wire2076 = {4'd3, 4'd2};
    assign wire2077 = {4'd3, 4'd2};
    assign wire2078 = {4'd3, 4'd2};
    assign wire2079 = {4'd3, 4'd2};
    assign wire2080 = {4'd4, 4'd2};
    assign wire2081 = {4'd4, 4'd2};
    assign wire2082 = {4'd4, 4'd2};
    assign wire2083 = {4'd4, 4'd2};
    assign wire2084 = {4'd4, 4'd2};
    assign wire2085 = {4'd4, 4'd2};
    assign wire2086 = {4'd4, 4'd2};
    assign wire2087 = {4'd4, 4'd2};
    assign wire2088 = {4'd4, 4'd2};
    assign wire2089 = {4'd4, 4'd2};
    assign wire2090 = {4'd4, 4'd2};
    assign wire2091 = {4'd4, 4'd2};
    assign wire2092 = {4'd4, 4'd2};
    assign wire2093 = {4'd4, 4'd2};
    assign wire2094 = {4'd4, 4'd2};
    assign wire2095 = {4'd4, 4'd2};
    assign wire2096 = {4'd4, 4'd2};
    assign wire2097 = {4'd4, 4'd2};
    assign wire2098 = {4'd4, 4'd2};
    assign wire2099 = {4'd4, 4'd2};
    assign wire2100 = {4'd4, 4'd2};
    assign wire2101 = {4'd4, 4'd2};
    assign wire2102 = {4'd4, 4'd2};
    assign wire2103 = {4'd4, 4'd2};
    assign wire2104 = {4'd4, 4'd2};
    assign wire2105 = {4'd4, 4'd2};
    assign wire2106 = {4'd4, 4'd2};
    assign wire2107 = {4'd4, 4'd2};
    assign wire2108 = {4'd4, 4'd2};
    assign wire2109 = {4'd4, 4'd2};
    assign wire2110 = {4'd4, 4'd2};
    assign wire2111 = {4'd4, 4'd2};
    assign wire2112 = {4'd6, 4'd2};
    assign wire2113 = {4'd6, 4'd2};
    assign wire2114 = {4'd6, 4'd2};
    assign wire2115 = {4'd6, 4'd2};
    assign wire2116 = {4'd6, 4'd2};
    assign wire2117 = {4'd6, 4'd2};
    assign wire2118 = {4'd6, 4'd2};
    assign wire2119 = {4'd6, 4'd2};
    assign wire2120 = {4'd6, 4'd2};
    assign wire2121 = {4'd6, 4'd2};
    assign wire2122 = {4'd6, 4'd2};
    assign wire2123 = {4'd6, 4'd2};
    assign wire2124 = {4'd6, 4'd2};
    assign wire2125 = {4'd6, 4'd2};
    assign wire2126 = {4'd6, 4'd2};
    assign wire2127 = {4'd6, 4'd2};
    assign wire2128 = {4'd6, 4'd2};
    assign wire2129 = {4'd6, 4'd2};
    assign wire2130 = {4'd6, 4'd2};
    assign wire2131 = {4'd6, 4'd2};
    assign wire2132 = {4'd6, 4'd2};
    assign wire2133 = {4'd6, 4'd2};
    assign wire2134 = {4'd6, 4'd2};
    assign wire2135 = {4'd6, 4'd2};
    assign wire2136 = {4'd6, 4'd2};
    assign wire2137 = {4'd6, 4'd2};
    assign wire2138 = {4'd6, 4'd2};
    assign wire2139 = {4'd6, 4'd2};
    assign wire2140 = {4'd6, 4'd2};
    assign wire2141 = {4'd6, 4'd2};
    assign wire2142 = {4'd6, 4'd2};
    assign wire2143 = {4'd6, 4'd2};
    assign wire2144 = {4'd8, 4'd2};
    assign wire2145 = {4'd8, 4'd2};
    assign wire2146 = {4'd8, 4'd2};
    assign wire2147 = {4'd8, 4'd2};
    assign wire2148 = {4'd8, 4'd2};
    assign wire2149 = {4'd8, 4'd2};
    assign wire2150 = {4'd8, 4'd2};
    assign wire2151 = {4'd8, 4'd2};
    assign wire2152 = {4'd8, 4'd2};
    assign wire2153 = {4'd8, 4'd2};
    assign wire2154 = {4'd8, 4'd2};
    assign wire2155 = {4'd8, 4'd2};
    assign wire2156 = {4'd8, 4'd2};
    assign wire2157 = {4'd8, 4'd2};
    assign wire2158 = {4'd8, 4'd2};
    assign wire2159 = {4'd8, 4'd2};
    assign wire2160 = {4'd8, 4'd2};
    assign wire2161 = {4'd8, 4'd2};
    assign wire2162 = {4'd8, 4'd2};
    assign wire2163 = {4'd8, 4'd2};
    assign wire2164 = {4'd8, 4'd2};
    assign wire2165 = {4'd8, 4'd2};
    assign wire2166 = {4'd8, 4'd2};
    assign wire2167 = {4'd8, 4'd2};
    assign wire2168 = {4'd8, 4'd2};
    assign wire2169 = {4'd8, 4'd2};
    assign wire2170 = {4'd8, 4'd2};
    assign wire2171 = {4'd8, 4'd2};
    assign wire2172 = {4'd8, 4'd2};
    assign wire2173 = {4'd8, 4'd2};
    assign wire2174 = {4'd8, 4'd2};
    assign wire2175 = {4'd8, 4'd2};
    assign wire2176 = {4'd4, 4'd3};
    assign wire2177 = {4'd4, 4'd3};
    assign wire2178 = {4'd4, 4'd3};
    assign wire2179 = {4'd4, 4'd3};
    assign wire2180 = {4'd5, 4'd4};
    assign wire2181 = {4'd8, 4'd7};
    assign wire2182 = {4'd4, 4'd3};
    assign wire2183 = {4'd4, 4'd3};
    assign wire2184 = {4'd5, 4'd4};
    assign wire2185 = {4'd5, 4'd4};
    assign wire2186 = {4'd5, 4'd4};
    assign wire2187 = {4'd5, 4'd4};
    assign wire2188 = {4'd6, 4'd5};
    assign wire2189 = {4'd5, 4'd4};
    assign wire2190 = {4'd5, 4'd4};
    assign wire2191 = {4'd5, 4'd4};
    assign wire2192 = {4'd8, 4'd7};
    assign wire2193 = {4'd8, 4'd7};
    assign wire2194 = {4'd8, 4'd7};
    assign wire2195 = {4'd8, 4'd7};
    assign wire2196 = {4'd9, 4'd8};
    assign wire2197 = {4'd8, 4'd7};
    assign wire2198 = {4'd8, 4'd7};
    assign wire2199 = {4'd8, 4'd7};
    assign wire2200 = {4'd4, 4'd3};
    assign wire2201 = {4'd4, 4'd3};
    assign wire2202 = {4'd4, 4'd3};
    assign wire2203 = {4'd4, 4'd3};
    assign wire2204 = {4'd4, 4'd3};
    assign wire2205 = {4'd4, 4'd3};
    assign wire2206 = {4'd4, 4'd3};
    assign wire2207 = {4'd4, 4'd3};
    assign wire2208 = {4'd5, 4'd3};
    assign wire2209 = {4'd5, 4'd3};
    assign wire2210 = {4'd5, 4'd3};
    assign wire2211 = {4'd5, 4'd3};
    assign wire2212 = {4'd6, 4'd4};
    assign wire2213 = {4'd9, 4'd7};
    assign wire2214 = {4'd5, 4'd3};
    assign wire2215 = {4'd5, 4'd3};
    assign wire2216 = {4'd6, 4'd4};
    assign wire2217 = {4'd6, 4'd4};
    assign wire2218 = {4'd6, 4'd4};
    assign wire2219 = {4'd6, 4'd4};
    assign wire2220 = {4'd7, 4'd5};
    assign wire2221 = {4'd6, 4'd4};
    assign wire2222 = {4'd6, 4'd4};
    assign wire2223 = {4'd6, 4'd4};
    assign wire2224 = {4'd9, 4'd7};
    assign wire2225 = {4'd9, 4'd7};
    assign wire2226 = {4'd9, 4'd7};
    assign wire2227 = {4'd9, 4'd7};
    assign wire2228 = {4'd10, 4'd8};
    assign wire2229 = {4'd9, 4'd7};
    assign wire2230 = {4'd9, 4'd7};
    assign wire2231 = {4'd9, 4'd7};
    assign wire2232 = {4'd5, 4'd3};
    assign wire2233 = {4'd5, 4'd3};
    assign wire2234 = {4'd5, 4'd3};
    assign wire2235 = {4'd5, 4'd3};
    assign wire2236 = {4'd5, 4'd3};
    assign wire2237 = {4'd5, 4'd3};
    assign wire2238 = {4'd5, 4'd3};
    assign wire2239 = {4'd5, 4'd3};
    assign wire2240 = {4'd7, 4'd3};
    assign wire2241 = {4'd7, 4'd3};
    assign wire2242 = {4'd7, 4'd3};
    assign wire2243 = {4'd7, 4'd3};
    assign wire2244 = {4'd8, 4'd4};
    assign wire2245 = {4'd11, 4'd7};
    assign wire2246 = {4'd7, 4'd3};
    assign wire2247 = {4'd7, 4'd3};
    assign wire2248 = {4'd8, 4'd4};
    assign wire2249 = {4'd8, 4'd4};
    assign wire2250 = {4'd8, 4'd4};
    assign wire2251 = {4'd8, 4'd4};
    assign wire2252 = {4'd9, 4'd5};
    assign wire2253 = {4'd8, 4'd4};
    assign wire2254 = {4'd8, 4'd4};
    assign wire2255 = {4'd8, 4'd4};
    assign wire2256 = {4'd11, 4'd7};
    assign wire2257 = {4'd11, 4'd7};
    assign wire2258 = {4'd11, 4'd7};
    assign wire2259 = {4'd11, 4'd7};
    assign wire2260 = {4'd12, 4'd8};
    assign wire2261 = {4'd11, 4'd7};
    assign wire2262 = {4'd11, 4'd7};
    assign wire2263 = {4'd11, 4'd7};
    assign wire2264 = {4'd7, 4'd3};
    assign wire2265 = {4'd7, 4'd3};
    assign wire2266 = {4'd7, 4'd3};
    assign wire2267 = {4'd7, 4'd3};
    assign wire2268 = {4'd7, 4'd3};
    assign wire2269 = {4'd7, 4'd3};
    assign wire2270 = {4'd7, 4'd3};
    assign wire2271 = {4'd7, 4'd3};
    assign wire2272 = {4'd9, 4'd3};
    assign wire2273 = {4'd9, 4'd3};
    assign wire2274 = {4'd9, 4'd3};
    assign wire2275 = {4'd9, 4'd3};
    assign wire2276 = {4'd10, 4'd4};
    assign wire2277 = {4'd13, 4'd7};
    assign wire2278 = {4'd9, 4'd3};
    assign wire2279 = {4'd9, 4'd3};
    assign wire2280 = {4'd10, 4'd4};
    assign wire2281 = {4'd10, 4'd4};
    assign wire2282 = {4'd10, 4'd4};
    assign wire2283 = {4'd10, 4'd4};
    assign wire2284 = {4'd11, 4'd5};
    assign wire2285 = {4'd10, 4'd4};
    assign wire2286 = {4'd10, 4'd4};
    assign wire2287 = {4'd10, 4'd4};
    assign wire2288 = {4'd13, 4'd7};
    assign wire2289 = {4'd13, 4'd7};
    assign wire2290 = {4'd13, 4'd7};
    assign wire2291 = {4'd13, 4'd7};
    assign wire2292 = {4'd14, 4'd8};
    assign wire2293 = {4'd13, 4'd7};
    assign wire2294 = {4'd13, 4'd7};
    assign wire2295 = {4'd13, 4'd7};
    assign wire2296 = {4'd9, 4'd3};
    assign wire2297 = {4'd9, 4'd3};
    assign wire2298 = {4'd9, 4'd3};
    assign wire2299 = {4'd9, 4'd3};
    assign wire2300 = {4'd9, 4'd3};
    assign wire2301 = {4'd9, 4'd3};
    assign wire2302 = {4'd9, 4'd3};
    assign wire2303 = {4'd9, 4'd3};
    assign wire2304 = {4'd4, 4'd3};
    assign wire2305 = {4'd4, 4'd3};
    assign wire2306 = {4'd4, 4'd3};
    assign wire2307 = {4'd4, 4'd3};
    assign wire2308 = {4'd4, 4'd3};
    assign wire2309 = {4'd4, 4'd3};
    assign wire2310 = {4'd4, 4'd3};
    assign wire2311 = {4'd4, 4'd3};
    assign wire2312 = {4'd4, 4'd3};
    assign wire2313 = {4'd4, 4'd3};
    assign wire2314 = {4'd4, 4'd3};
    assign wire2315 = {4'd4, 4'd3};
    assign wire2316 = {4'd4, 4'd3};
    assign wire2317 = {4'd4, 4'd3};
    assign wire2318 = {4'd4, 4'd3};
    assign wire2319 = {4'd4, 4'd3};
    assign wire2320 = {4'd4, 4'd3};
    assign wire2321 = {4'd4, 4'd3};
    assign wire2322 = {4'd4, 4'd3};
    assign wire2323 = {4'd4, 4'd3};
    assign wire2324 = {4'd4, 4'd3};
    assign wire2325 = {4'd4, 4'd3};
    assign wire2326 = {4'd4, 4'd3};
    assign wire2327 = {4'd4, 4'd3};
    assign wire2328 = {4'd4, 4'd3};
    assign wire2329 = {4'd4, 4'd3};
    assign wire2330 = {4'd4, 4'd3};
    assign wire2331 = {4'd4, 4'd3};
    assign wire2332 = {4'd4, 4'd3};
    assign wire2333 = {4'd4, 4'd3};
    assign wire2334 = {4'd4, 4'd3};
    assign wire2335 = {4'd4, 4'd3};
    assign wire2336 = {4'd5, 4'd3};
    assign wire2337 = {4'd5, 4'd3};
    assign wire2338 = {4'd5, 4'd3};
    assign wire2339 = {4'd5, 4'd3};
    assign wire2340 = {4'd5, 4'd3};
    assign wire2341 = {4'd5, 4'd3};
    assign wire2342 = {4'd5, 4'd3};
    assign wire2343 = {4'd5, 4'd3};
    assign wire2344 = {4'd5, 4'd3};
    assign wire2345 = {4'd5, 4'd3};
    assign wire2346 = {4'd5, 4'd3};
    assign wire2347 = {4'd5, 4'd3};
    assign wire2348 = {4'd5, 4'd3};
    assign wire2349 = {4'd5, 4'd3};
    assign wire2350 = {4'd5, 4'd3};
    assign wire2351 = {4'd5, 4'd3};
    assign wire2352 = {4'd5, 4'd3};
    assign wire2353 = {4'd5, 4'd3};
    assign wire2354 = {4'd5, 4'd3};
    assign wire2355 = {4'd5, 4'd3};
    assign wire2356 = {4'd5, 4'd3};
    assign wire2357 = {4'd5, 4'd3};
    assign wire2358 = {4'd5, 4'd3};
    assign wire2359 = {4'd5, 4'd3};
    assign wire2360 = {4'd5, 4'd3};
    assign wire2361 = {4'd5, 4'd3};
    assign wire2362 = {4'd5, 4'd3};
    assign wire2363 = {4'd5, 4'd3};
    assign wire2364 = {4'd5, 4'd3};
    assign wire2365 = {4'd5, 4'd3};
    assign wire2366 = {4'd5, 4'd3};
    assign wire2367 = {4'd5, 4'd3};
    assign wire2368 = {4'd7, 4'd3};
    assign wire2369 = {4'd7, 4'd3};
    assign wire2370 = {4'd7, 4'd3};
    assign wire2371 = {4'd7, 4'd3};
    assign wire2372 = {4'd7, 4'd3};
    assign wire2373 = {4'd7, 4'd3};
    assign wire2374 = {4'd7, 4'd3};
    assign wire2375 = {4'd7, 4'd3};
    assign wire2376 = {4'd7, 4'd3};
    assign wire2377 = {4'd7, 4'd3};
    assign wire2378 = {4'd7, 4'd3};
    assign wire2379 = {4'd7, 4'd3};
    assign wire2380 = {4'd7, 4'd3};
    assign wire2381 = {4'd7, 4'd3};
    assign wire2382 = {4'd7, 4'd3};
    assign wire2383 = {4'd7, 4'd3};
    assign wire2384 = {4'd7, 4'd3};
    assign wire2385 = {4'd7, 4'd3};
    assign wire2386 = {4'd7, 4'd3};
    assign wire2387 = {4'd7, 4'd3};
    assign wire2388 = {4'd7, 4'd3};
    assign wire2389 = {4'd7, 4'd3};
    assign wire2390 = {4'd7, 4'd3};
    assign wire2391 = {4'd7, 4'd3};
    assign wire2392 = {4'd7, 4'd3};
    assign wire2393 = {4'd7, 4'd3};
    assign wire2394 = {4'd7, 4'd3};
    assign wire2395 = {4'd7, 4'd3};
    assign wire2396 = {4'd7, 4'd3};
    assign wire2397 = {4'd7, 4'd3};
    assign wire2398 = {4'd7, 4'd3};
    assign wire2399 = {4'd7, 4'd3};
    assign wire2400 = {4'd9, 4'd3};
    assign wire2401 = {4'd9, 4'd3};
    assign wire2402 = {4'd9, 4'd3};
    assign wire2403 = {4'd9, 4'd3};
    assign wire2404 = {4'd9, 4'd3};
    assign wire2405 = {4'd9, 4'd3};
    assign wire2406 = {4'd9, 4'd3};
    assign wire2407 = {4'd9, 4'd3};
    assign wire2408 = {4'd9, 4'd3};
    assign wire2409 = {4'd9, 4'd3};
    assign wire2410 = {4'd9, 4'd3};
    assign wire2411 = {4'd9, 4'd3};
    assign wire2412 = {4'd9, 4'd3};
    assign wire2413 = {4'd9, 4'd3};
    assign wire2414 = {4'd9, 4'd3};
    assign wire2415 = {4'd9, 4'd3};
    assign wire2416 = {4'd9, 4'd3};
    assign wire2417 = {4'd9, 4'd3};
    assign wire2418 = {4'd9, 4'd3};
    assign wire2419 = {4'd9, 4'd3};
    assign wire2420 = {4'd9, 4'd3};
    assign wire2421 = {4'd9, 4'd3};
    assign wire2422 = {4'd9, 4'd3};
    assign wire2423 = {4'd9, 4'd3};
    assign wire2424 = {4'd9, 4'd3};
    assign wire2425 = {4'd9, 4'd3};
    assign wire2426 = {4'd9, 4'd3};
    assign wire2427 = {4'd9, 4'd3};
    assign wire2428 = {4'd9, 4'd3};
    assign wire2429 = {4'd9, 4'd3};
    assign wire2430 = {4'd9, 4'd3};
    assign wire2431 = {4'd9, 4'd3};
    assign wire2432 = {4'd5, 4'd4};
    assign wire2433 = {4'd5, 4'd4};
    assign wire2434 = {4'd5, 4'd4};
    assign wire2435 = {4'd5, 4'd4};
    assign wire2436 = {4'd6, 4'd5};
    assign wire2437 = {4'd9, 4'd8};
    assign wire2438 = {4'd5, 4'd4};
    assign wire2439 = {4'd5, 4'd4};
    assign wire2440 = {4'd6, 4'd5};
    assign wire2441 = {4'd6, 4'd5};
    assign wire2442 = {4'd6, 4'd5};
    assign wire2443 = {4'd6, 4'd5};
    assign wire2444 = {4'd7, 4'd6};
    assign wire2445 = {4'd6, 4'd5};
    assign wire2446 = {4'd6, 4'd5};
    assign wire2447 = {4'd6, 4'd5};
    assign wire2448 = {4'd9, 4'd8};
    assign wire2449 = {4'd9, 4'd8};
    assign wire2450 = {4'd9, 4'd8};
    assign wire2451 = {4'd9, 4'd8};
    assign wire2452 = {4'd10, 4'd9};
    assign wire2453 = {4'd9, 4'd8};
    assign wire2454 = {4'd9, 4'd8};
    assign wire2455 = {4'd9, 4'd8};
    assign wire2456 = {4'd5, 4'd4};
    assign wire2457 = {4'd5, 4'd4};
    assign wire2458 = {4'd5, 4'd4};
    assign wire2459 = {4'd5, 4'd4};
    assign wire2460 = {4'd5, 4'd4};
    assign wire2461 = {4'd5, 4'd4};
    assign wire2462 = {4'd5, 4'd4};
    assign wire2463 = {4'd5, 4'd4};
    assign wire2464 = {4'd6, 4'd4};
    assign wire2465 = {4'd6, 4'd4};
    assign wire2466 = {4'd6, 4'd4};
    assign wire2467 = {4'd6, 4'd4};
    assign wire2468 = {4'd7, 4'd5};
    assign wire2469 = {4'd10, 4'd8};
    assign wire2470 = {4'd6, 4'd4};
    assign wire2471 = {4'd6, 4'd4};
    assign wire2472 = {4'd7, 4'd5};
    assign wire2473 = {4'd7, 4'd5};
    assign wire2474 = {4'd7, 4'd5};
    assign wire2475 = {4'd7, 4'd5};
    assign wire2476 = {4'd8, 4'd6};
    assign wire2477 = {4'd7, 4'd5};
    assign wire2478 = {4'd7, 4'd5};
    assign wire2479 = {4'd7, 4'd5};
    assign wire2480 = {4'd10, 4'd8};
    assign wire2481 = {4'd10, 4'd8};
    assign wire2482 = {4'd10, 4'd8};
    assign wire2483 = {4'd10, 4'd8};
    assign wire2484 = {4'd11, 4'd9};
    assign wire2485 = {4'd10, 4'd8};
    assign wire2486 = {4'd10, 4'd8};
    assign wire2487 = {4'd10, 4'd8};
    assign wire2488 = {4'd6, 4'd4};
    assign wire2489 = {4'd6, 4'd4};
    assign wire2490 = {4'd6, 4'd4};
    assign wire2491 = {4'd6, 4'd4};
    assign wire2492 = {4'd6, 4'd4};
    assign wire2493 = {4'd6, 4'd4};
    assign wire2494 = {4'd6, 4'd4};
    assign wire2495 = {4'd6, 4'd4};
    assign wire2496 = {4'd8, 4'd4};
    assign wire2497 = {4'd8, 4'd4};
    assign wire2498 = {4'd8, 4'd4};
    assign wire2499 = {4'd8, 4'd4};
    assign wire2500 = {4'd9, 4'd5};
    assign wire2501 = {4'd12, 4'd8};
    assign wire2502 = {4'd8, 4'd4};
    assign wire2503 = {4'd8, 4'd4};
    assign wire2504 = {4'd9, 4'd5};
    assign wire2505 = {4'd9, 4'd5};
    assign wire2506 = {4'd9, 4'd5};
    assign wire2507 = {4'd9, 4'd5};
    assign wire2508 = {4'd10, 4'd6};
    assign wire2509 = {4'd9, 4'd5};
    assign wire2510 = {4'd9, 4'd5};
    assign wire2511 = {4'd9, 4'd5};
    assign wire2512 = {4'd12, 4'd8};
    assign wire2513 = {4'd12, 4'd8};
    assign wire2514 = {4'd12, 4'd8};
    assign wire2515 = {4'd12, 4'd8};
    assign wire2516 = {4'd13, 4'd9};
    assign wire2517 = {4'd12, 4'd8};
    assign wire2518 = {4'd12, 4'd8};
    assign wire2519 = {4'd12, 4'd8};
    assign wire2520 = {4'd8, 4'd4};
    assign wire2521 = {4'd8, 4'd4};
    assign wire2522 = {4'd8, 4'd4};
    assign wire2523 = {4'd8, 4'd4};
    assign wire2524 = {4'd8, 4'd4};
    assign wire2525 = {4'd8, 4'd4};
    assign wire2526 = {4'd8, 4'd4};
    assign wire2527 = {4'd8, 4'd4};
    assign wire2528 = {4'd10, 4'd4};
    assign wire2529 = {4'd10, 4'd4};
    assign wire2530 = {4'd10, 4'd4};
    assign wire2531 = {4'd10, 4'd4};
    assign wire2532 = {4'd11, 4'd5};
    assign wire2533 = {4'd14, 4'd8};
    assign wire2534 = {4'd10, 4'd4};
    assign wire2535 = {4'd10, 4'd4};
    assign wire2536 = {4'd11, 4'd5};
    assign wire2537 = {4'd11, 4'd5};
    assign wire2538 = {4'd11, 4'd5};
    assign wire2539 = {4'd11, 4'd5};
    assign wire2540 = {4'd12, 4'd6};
    assign wire2541 = {4'd11, 4'd5};
    assign wire2542 = {4'd11, 4'd5};
    assign wire2543 = {4'd11, 4'd5};
    assign wire2544 = {4'd14, 4'd8};
    assign wire2545 = {4'd14, 4'd8};
    assign wire2546 = {4'd14, 4'd8};
    assign wire2547 = {4'd14, 4'd8};
    assign wire2548 = {4'd15, 4'd9};
    assign wire2549 = {4'd14, 4'd8};
    assign wire2550 = {4'd14, 4'd8};
    assign wire2551 = {4'd14, 4'd8};
    assign wire2552 = {4'd10, 4'd4};
    assign wire2553 = {4'd10, 4'd4};
    assign wire2554 = {4'd10, 4'd4};
    assign wire2555 = {4'd10, 4'd4};
    assign wire2556 = {4'd10, 4'd4};
    assign wire2557 = {4'd10, 4'd4};
    assign wire2558 = {4'd10, 4'd4};
    assign wire2559 = {4'd10, 4'd4};
    assign wire2560 = {4'd4, 4'd3};
    assign wire2561 = {4'd4, 4'd3};
    assign wire2562 = {4'd4, 4'd3};
    assign wire2563 = {4'd4, 4'd3};
    assign wire2564 = {4'd4, 4'd3};
    assign wire2565 = {4'd4, 4'd3};
    assign wire2566 = {4'd4, 4'd3};
    assign wire2567 = {4'd4, 4'd3};
    assign wire2568 = {4'd4, 4'd3};
    assign wire2569 = {4'd4, 4'd3};
    assign wire2570 = {4'd4, 4'd3};
    assign wire2571 = {4'd4, 4'd3};
    assign wire2572 = {4'd4, 4'd3};
    assign wire2573 = {4'd4, 4'd3};
    assign wire2574 = {4'd4, 4'd3};
    assign wire2575 = {4'd4, 4'd3};
    assign wire2576 = {4'd4, 4'd3};
    assign wire2577 = {4'd4, 4'd3};
    assign wire2578 = {4'd4, 4'd3};
    assign wire2579 = {4'd4, 4'd3};
    assign wire2580 = {4'd4, 4'd3};
    assign wire2581 = {4'd4, 4'd3};
    assign wire2582 = {4'd4, 4'd3};
    assign wire2583 = {4'd4, 4'd3};
    assign wire2584 = {4'd4, 4'd3};
    assign wire2585 = {4'd4, 4'd3};
    assign wire2586 = {4'd4, 4'd3};
    assign wire2587 = {4'd4, 4'd3};
    assign wire2588 = {4'd4, 4'd3};
    assign wire2589 = {4'd4, 4'd3};
    assign wire2590 = {4'd4, 4'd3};
    assign wire2591 = {4'd4, 4'd3};
    assign wire2592 = {4'd5, 4'd3};
    assign wire2593 = {4'd5, 4'd3};
    assign wire2594 = {4'd5, 4'd3};
    assign wire2595 = {4'd5, 4'd3};
    assign wire2596 = {4'd5, 4'd3};
    assign wire2597 = {4'd5, 4'd3};
    assign wire2598 = {4'd5, 4'd3};
    assign wire2599 = {4'd5, 4'd3};
    assign wire2600 = {4'd5, 4'd3};
    assign wire2601 = {4'd5, 4'd3};
    assign wire2602 = {4'd5, 4'd3};
    assign wire2603 = {4'd5, 4'd3};
    assign wire2604 = {4'd5, 4'd3};
    assign wire2605 = {4'd5, 4'd3};
    assign wire2606 = {4'd5, 4'd3};
    assign wire2607 = {4'd5, 4'd3};
    assign wire2608 = {4'd5, 4'd3};
    assign wire2609 = {4'd5, 4'd3};
    assign wire2610 = {4'd5, 4'd3};
    assign wire2611 = {4'd5, 4'd3};
    assign wire2612 = {4'd5, 4'd3};
    assign wire2613 = {4'd5, 4'd3};
    assign wire2614 = {4'd5, 4'd3};
    assign wire2615 = {4'd5, 4'd3};
    assign wire2616 = {4'd5, 4'd3};
    assign wire2617 = {4'd5, 4'd3};
    assign wire2618 = {4'd5, 4'd3};
    assign wire2619 = {4'd5, 4'd3};
    assign wire2620 = {4'd5, 4'd3};
    assign wire2621 = {4'd5, 4'd3};
    assign wire2622 = {4'd5, 4'd3};
    assign wire2623 = {4'd5, 4'd3};
    assign wire2624 = {4'd7, 4'd3};
    assign wire2625 = {4'd7, 4'd3};
    assign wire2626 = {4'd7, 4'd3};
    assign wire2627 = {4'd7, 4'd3};
    assign wire2628 = {4'd7, 4'd3};
    assign wire2629 = {4'd7, 4'd3};
    assign wire2630 = {4'd7, 4'd3};
    assign wire2631 = {4'd7, 4'd3};
    assign wire2632 = {4'd7, 4'd3};
    assign wire2633 = {4'd7, 4'd3};
    assign wire2634 = {4'd7, 4'd3};
    assign wire2635 = {4'd7, 4'd3};
    assign wire2636 = {4'd7, 4'd3};
    assign wire2637 = {4'd7, 4'd3};
    assign wire2638 = {4'd7, 4'd3};
    assign wire2639 = {4'd7, 4'd3};
    assign wire2640 = {4'd7, 4'd3};
    assign wire2641 = {4'd7, 4'd3};
    assign wire2642 = {4'd7, 4'd3};
    assign wire2643 = {4'd7, 4'd3};
    assign wire2644 = {4'd7, 4'd3};
    assign wire2645 = {4'd7, 4'd3};
    assign wire2646 = {4'd7, 4'd3};
    assign wire2647 = {4'd7, 4'd3};
    assign wire2648 = {4'd7, 4'd3};
    assign wire2649 = {4'd7, 4'd3};
    assign wire2650 = {4'd7, 4'd3};
    assign wire2651 = {4'd7, 4'd3};
    assign wire2652 = {4'd7, 4'd3};
    assign wire2653 = {4'd7, 4'd3};
    assign wire2654 = {4'd7, 4'd3};
    assign wire2655 = {4'd7, 4'd3};
    assign wire2656 = {4'd9, 4'd3};
    assign wire2657 = {4'd9, 4'd3};
    assign wire2658 = {4'd9, 4'd3};
    assign wire2659 = {4'd9, 4'd3};
    assign wire2660 = {4'd9, 4'd3};
    assign wire2661 = {4'd9, 4'd3};
    assign wire2662 = {4'd9, 4'd3};
    assign wire2663 = {4'd9, 4'd3};
    assign wire2664 = {4'd9, 4'd3};
    assign wire2665 = {4'd9, 4'd3};
    assign wire2666 = {4'd9, 4'd3};
    assign wire2667 = {4'd9, 4'd3};
    assign wire2668 = {4'd9, 4'd3};
    assign wire2669 = {4'd9, 4'd3};
    assign wire2670 = {4'd9, 4'd3};
    assign wire2671 = {4'd9, 4'd3};
    assign wire2672 = {4'd9, 4'd3};
    assign wire2673 = {4'd9, 4'd3};
    assign wire2674 = {4'd9, 4'd3};
    assign wire2675 = {4'd9, 4'd3};
    assign wire2676 = {4'd9, 4'd3};
    assign wire2677 = {4'd9, 4'd3};
    assign wire2678 = {4'd9, 4'd3};
    assign wire2679 = {4'd9, 4'd3};
    assign wire2680 = {4'd9, 4'd3};
    assign wire2681 = {4'd9, 4'd3};
    assign wire2682 = {4'd9, 4'd3};
    assign wire2683 = {4'd9, 4'd3};
    assign wire2684 = {4'd9, 4'd3};
    assign wire2685 = {4'd9, 4'd3};
    assign wire2686 = {4'd9, 4'd3};
    assign wire2687 = {4'd9, 4'd3};
    assign wire2688 = {4'd5, 4'd4};
    assign wire2689 = {4'd5, 4'd4};
    assign wire2690 = {4'd5, 4'd4};
    assign wire2691 = {4'd5, 4'd4};
    assign wire2692 = {4'd5, 4'd4};
    assign wire2693 = {4'd7, 4'd6};
    assign wire2694 = {4'd5, 4'd4};
    assign wire2695 = {4'd5, 4'd4};
    assign wire2696 = {4'd6, 4'd5};
    assign wire2697 = {4'd6, 4'd5};
    assign wire2698 = {4'd6, 4'd5};
    assign wire2699 = {4'd6, 4'd5};
    assign wire2700 = {4'd6, 4'd5};
    assign wire2701 = {4'd6, 4'd5};
    assign wire2702 = {4'd6, 4'd5};
    assign wire2703 = {4'd6, 4'd5};
    assign wire2704 = {4'd7, 4'd6};
    assign wire2705 = {4'd7, 4'd6};
    assign wire2706 = {4'd7, 4'd6};
    assign wire2707 = {4'd7, 4'd6};
    assign wire2708 = {4'd7, 4'd6};
    assign wire2709 = {4'd7, 4'd6};
    assign wire2710 = {4'd7, 4'd6};
    assign wire2711 = {4'd7, 4'd6};
    assign wire2712 = {4'd5, 4'd4};
    assign wire2713 = {4'd5, 4'd4};
    assign wire2714 = {4'd5, 4'd4};
    assign wire2715 = {4'd5, 4'd4};
    assign wire2716 = {4'd5, 4'd4};
    assign wire2717 = {4'd5, 4'd4};
    assign wire2718 = {4'd5, 4'd4};
    assign wire2719 = {4'd5, 4'd4};
    assign wire2720 = {4'd6, 4'd4};
    assign wire2721 = {4'd6, 4'd4};
    assign wire2722 = {4'd6, 4'd4};
    assign wire2723 = {4'd6, 4'd4};
    assign wire2724 = {4'd6, 4'd4};
    assign wire2725 = {4'd8, 4'd6};
    assign wire2726 = {4'd6, 4'd4};
    assign wire2727 = {4'd6, 4'd4};
    assign wire2728 = {4'd7, 4'd5};
    assign wire2729 = {4'd7, 4'd5};
    assign wire2730 = {4'd7, 4'd5};
    assign wire2731 = {4'd7, 4'd5};
    assign wire2732 = {4'd7, 4'd5};
    assign wire2733 = {4'd7, 4'd5};
    assign wire2734 = {4'd7, 4'd5};
    assign wire2735 = {4'd7, 4'd5};
    assign wire2736 = {4'd8, 4'd6};
    assign wire2737 = {4'd8, 4'd6};
    assign wire2738 = {4'd8, 4'd6};
    assign wire2739 = {4'd8, 4'd6};
    assign wire2740 = {4'd8, 4'd6};
    assign wire2741 = {4'd8, 4'd6};
    assign wire2742 = {4'd8, 4'd6};
    assign wire2743 = {4'd8, 4'd6};
    assign wire2744 = {4'd6, 4'd4};
    assign wire2745 = {4'd6, 4'd4};
    assign wire2746 = {4'd6, 4'd4};
    assign wire2747 = {4'd6, 4'd4};
    assign wire2748 = {4'd6, 4'd4};
    assign wire2749 = {4'd6, 4'd4};
    assign wire2750 = {4'd6, 4'd4};
    assign wire2751 = {4'd6, 4'd4};
    assign wire2752 = {4'd8, 4'd4};
    assign wire2753 = {4'd8, 4'd4};
    assign wire2754 = {4'd8, 4'd4};
    assign wire2755 = {4'd8, 4'd4};
    assign wire2756 = {4'd8, 4'd4};
    assign wire2757 = {4'd10, 4'd6};
    assign wire2758 = {4'd8, 4'd4};
    assign wire2759 = {4'd8, 4'd4};
    assign wire2760 = {4'd9, 4'd5};
    assign wire2761 = {4'd9, 4'd5};
    assign wire2762 = {4'd9, 4'd5};
    assign wire2763 = {4'd9, 4'd5};
    assign wire2764 = {4'd9, 4'd5};
    assign wire2765 = {4'd9, 4'd5};
    assign wire2766 = {4'd9, 4'd5};
    assign wire2767 = {4'd9, 4'd5};
    assign wire2768 = {4'd10, 4'd6};
    assign wire2769 = {4'd10, 4'd6};
    assign wire2770 = {4'd10, 4'd6};
    assign wire2771 = {4'd10, 4'd6};
    assign wire2772 = {4'd10, 4'd6};
    assign wire2773 = {4'd10, 4'd6};
    assign wire2774 = {4'd10, 4'd6};
    assign wire2775 = {4'd10, 4'd6};
    assign wire2776 = {4'd8, 4'd4};
    assign wire2777 = {4'd8, 4'd4};
    assign wire2778 = {4'd8, 4'd4};
    assign wire2779 = {4'd8, 4'd4};
    assign wire2780 = {4'd8, 4'd4};
    assign wire2781 = {4'd8, 4'd4};
    assign wire2782 = {4'd8, 4'd4};
    assign wire2783 = {4'd8, 4'd4};
    assign wire2784 = {4'd10, 4'd4};
    assign wire2785 = {4'd10, 4'd4};
    assign wire2786 = {4'd10, 4'd4};
    assign wire2787 = {4'd10, 4'd4};
    assign wire2788 = {4'd10, 4'd4};
    assign wire2789 = {4'd12, 4'd6};
    assign wire2790 = {4'd10, 4'd4};
    assign wire2791 = {4'd10, 4'd4};
    assign wire2792 = {4'd11, 4'd5};
    assign wire2793 = {4'd11, 4'd5};
    assign wire2794 = {4'd11, 4'd5};
    assign wire2795 = {4'd11, 4'd5};
    assign wire2796 = {4'd11, 4'd5};
    assign wire2797 = {4'd11, 4'd5};
    assign wire2798 = {4'd11, 4'd5};
    assign wire2799 = {4'd11, 4'd5};
    assign wire2800 = {4'd12, 4'd6};
    assign wire2801 = {4'd12, 4'd6};
    assign wire2802 = {4'd12, 4'd6};
    assign wire2803 = {4'd12, 4'd6};
    assign wire2804 = {4'd12, 4'd6};
    assign wire2805 = {4'd12, 4'd6};
    assign wire2806 = {4'd12, 4'd6};
    assign wire2807 = {4'd12, 4'd6};
    assign wire2808 = {4'd10, 4'd4};
    assign wire2809 = {4'd10, 4'd4};
    assign wire2810 = {4'd10, 4'd4};
    assign wire2811 = {4'd10, 4'd4};
    assign wire2812 = {4'd10, 4'd4};
    assign wire2813 = {4'd10, 4'd4};
    assign wire2814 = {4'd10, 4'd4};
    assign wire2815 = {4'd10, 4'd4};
    assign wire2816 = {4'd5, 4'd4};
    assign wire2817 = {4'd5, 4'd4};
    assign wire2818 = {4'd5, 4'd4};
    assign wire2819 = {4'd5, 4'd4};
    assign wire2820 = {4'd5, 4'd4};
    assign wire2821 = {4'd5, 4'd4};
    assign wire2822 = {4'd5, 4'd4};
    assign wire2823 = {4'd5, 4'd4};
    assign wire2824 = {4'd5, 4'd4};
    assign wire2825 = {4'd5, 4'd4};
    assign wire2826 = {4'd5, 4'd4};
    assign wire2827 = {4'd5, 4'd4};
    assign wire2828 = {4'd5, 4'd4};
    assign wire2829 = {4'd5, 4'd4};
    assign wire2830 = {4'd5, 4'd4};
    assign wire2831 = {4'd5, 4'd4};
    assign wire2832 = {4'd5, 4'd4};
    assign wire2833 = {4'd5, 4'd4};
    assign wire2834 = {4'd5, 4'd4};
    assign wire2835 = {4'd5, 4'd4};
    assign wire2836 = {4'd5, 4'd4};
    assign wire2837 = {4'd5, 4'd4};
    assign wire2838 = {4'd5, 4'd4};
    assign wire2839 = {4'd5, 4'd4};
    assign wire2840 = {4'd5, 4'd4};
    assign wire2841 = {4'd5, 4'd4};
    assign wire2842 = {4'd5, 4'd4};
    assign wire2843 = {4'd5, 4'd4};
    assign wire2844 = {4'd5, 4'd4};
    assign wire2845 = {4'd5, 4'd4};
    assign wire2846 = {4'd5, 4'd4};
    assign wire2847 = {4'd5, 4'd4};
    assign wire2848 = {4'd6, 4'd4};
    assign wire2849 = {4'd6, 4'd4};
    assign wire2850 = {4'd6, 4'd4};
    assign wire2851 = {4'd6, 4'd4};
    assign wire2852 = {4'd6, 4'd4};
    assign wire2853 = {4'd6, 4'd4};
    assign wire2854 = {4'd6, 4'd4};
    assign wire2855 = {4'd6, 4'd4};
    assign wire2856 = {4'd6, 4'd4};
    assign wire2857 = {4'd6, 4'd4};
    assign wire2858 = {4'd6, 4'd4};
    assign wire2859 = {4'd6, 4'd4};
    assign wire2860 = {4'd6, 4'd4};
    assign wire2861 = {4'd6, 4'd4};
    assign wire2862 = {4'd6, 4'd4};
    assign wire2863 = {4'd6, 4'd4};
    assign wire2864 = {4'd6, 4'd4};
    assign wire2865 = {4'd6, 4'd4};
    assign wire2866 = {4'd6, 4'd4};
    assign wire2867 = {4'd6, 4'd4};
    assign wire2868 = {4'd6, 4'd4};
    assign wire2869 = {4'd6, 4'd4};
    assign wire2870 = {4'd6, 4'd4};
    assign wire2871 = {4'd6, 4'd4};
    assign wire2872 = {4'd6, 4'd4};
    assign wire2873 = {4'd6, 4'd4};
    assign wire2874 = {4'd6, 4'd4};
    assign wire2875 = {4'd6, 4'd4};
    assign wire2876 = {4'd6, 4'd4};
    assign wire2877 = {4'd6, 4'd4};
    assign wire2878 = {4'd6, 4'd4};
    assign wire2879 = {4'd6, 4'd4};
    assign wire2880 = {4'd8, 4'd4};
    assign wire2881 = {4'd8, 4'd4};
    assign wire2882 = {4'd8, 4'd4};
    assign wire2883 = {4'd8, 4'd4};
    assign wire2884 = {4'd8, 4'd4};
    assign wire2885 = {4'd8, 4'd4};
    assign wire2886 = {4'd8, 4'd4};
    assign wire2887 = {4'd8, 4'd4};
    assign wire2888 = {4'd8, 4'd4};
    assign wire2889 = {4'd8, 4'd4};
    assign wire2890 = {4'd8, 4'd4};
    assign wire2891 = {4'd8, 4'd4};
    assign wire2892 = {4'd8, 4'd4};
    assign wire2893 = {4'd8, 4'd4};
    assign wire2894 = {4'd8, 4'd4};
    assign wire2895 = {4'd8, 4'd4};
    assign wire2896 = {4'd8, 4'd4};
    assign wire2897 = {4'd8, 4'd4};
    assign wire2898 = {4'd8, 4'd4};
    assign wire2899 = {4'd8, 4'd4};
    assign wire2900 = {4'd8, 4'd4};
    assign wire2901 = {4'd8, 4'd4};
    assign wire2902 = {4'd8, 4'd4};
    assign wire2903 = {4'd8, 4'd4};
    assign wire2904 = {4'd8, 4'd4};
    assign wire2905 = {4'd8, 4'd4};
    assign wire2906 = {4'd8, 4'd4};
    assign wire2907 = {4'd8, 4'd4};
    assign wire2908 = {4'd8, 4'd4};
    assign wire2909 = {4'd8, 4'd4};
    assign wire2910 = {4'd8, 4'd4};
    assign wire2911 = {4'd8, 4'd4};
    assign wire2912 = {4'd10, 4'd4};
    assign wire2913 = {4'd10, 4'd4};
    assign wire2914 = {4'd10, 4'd4};
    assign wire2915 = {4'd10, 4'd4};
    assign wire2916 = {4'd10, 4'd4};
    assign wire2917 = {4'd10, 4'd4};
    assign wire2918 = {4'd10, 4'd4};
    assign wire2919 = {4'd10, 4'd4};
    assign wire2920 = {4'd10, 4'd4};
    assign wire2921 = {4'd10, 4'd4};
    assign wire2922 = {4'd10, 4'd4};
    assign wire2923 = {4'd10, 4'd4};
    assign wire2924 = {4'd10, 4'd4};
    assign wire2925 = {4'd10, 4'd4};
    assign wire2926 = {4'd10, 4'd4};
    assign wire2927 = {4'd10, 4'd4};
    assign wire2928 = {4'd10, 4'd4};
    assign wire2929 = {4'd10, 4'd4};
    assign wire2930 = {4'd10, 4'd4};
    assign wire2931 = {4'd10, 4'd4};
    assign wire2932 = {4'd10, 4'd4};
    assign wire2933 = {4'd10, 4'd4};
    assign wire2934 = {4'd10, 4'd4};
    assign wire2935 = {4'd10, 4'd4};
    assign wire2936 = {4'd10, 4'd4};
    assign wire2937 = {4'd10, 4'd4};
    assign wire2938 = {4'd10, 4'd4};
    assign wire2939 = {4'd10, 4'd4};
    assign wire2940 = {4'd10, 4'd4};
    assign wire2941 = {4'd10, 4'd4};
    assign wire2942 = {4'd10, 4'd4};
    assign wire2943 = {4'd10, 4'd4};
    assign wire2944 = {4'd6, 4'd5};
    assign wire2945 = {4'd6, 4'd5};
    assign wire2946 = {4'd6, 4'd5};
    assign wire2947 = {4'd6, 4'd5};
    assign wire2948 = {4'd6, 4'd5};
    assign wire2949 = {4'd8, 4'd7};
    assign wire2950 = {4'd6, 4'd5};
    assign wire2951 = {4'd6, 4'd5};
    assign wire2952 = {4'd7, 4'd6};
    assign wire2953 = {4'd7, 4'd6};
    assign wire2954 = {4'd7, 4'd6};
    assign wire2955 = {4'd7, 4'd6};
    assign wire2956 = {4'd7, 4'd6};
    assign wire2957 = {4'd7, 4'd6};
    assign wire2958 = {4'd7, 4'd6};
    assign wire2959 = {4'd7, 4'd6};
    assign wire2960 = {4'd8, 4'd7};
    assign wire2961 = {4'd8, 4'd7};
    assign wire2962 = {4'd8, 4'd7};
    assign wire2963 = {4'd8, 4'd7};
    assign wire2964 = {4'd8, 4'd7};
    assign wire2965 = {4'd8, 4'd7};
    assign wire2966 = {4'd8, 4'd7};
    assign wire2967 = {4'd8, 4'd7};
    assign wire2968 = {4'd6, 4'd5};
    assign wire2969 = {4'd6, 4'd5};
    assign wire2970 = {4'd6, 4'd5};
    assign wire2971 = {4'd6, 4'd5};
    assign wire2972 = {4'd6, 4'd5};
    assign wire2973 = {4'd6, 4'd5};
    assign wire2974 = {4'd6, 4'd5};
    assign wire2975 = {4'd6, 4'd5};
    assign wire2976 = {4'd7, 4'd5};
    assign wire2977 = {4'd7, 4'd5};
    assign wire2978 = {4'd7, 4'd5};
    assign wire2979 = {4'd7, 4'd5};
    assign wire2980 = {4'd7, 4'd5};
    assign wire2981 = {4'd9, 4'd7};
    assign wire2982 = {4'd7, 4'd5};
    assign wire2983 = {4'd7, 4'd5};
    assign wire2984 = {4'd8, 4'd6};
    assign wire2985 = {4'd8, 4'd6};
    assign wire2986 = {4'd8, 4'd6};
    assign wire2987 = {4'd8, 4'd6};
    assign wire2988 = {4'd8, 4'd6};
    assign wire2989 = {4'd8, 4'd6};
    assign wire2990 = {4'd8, 4'd6};
    assign wire2991 = {4'd8, 4'd6};
    assign wire2992 = {4'd9, 4'd7};
    assign wire2993 = {4'd9, 4'd7};
    assign wire2994 = {4'd9, 4'd7};
    assign wire2995 = {4'd9, 4'd7};
    assign wire2996 = {4'd9, 4'd7};
    assign wire2997 = {4'd9, 4'd7};
    assign wire2998 = {4'd9, 4'd7};
    assign wire2999 = {4'd9, 4'd7};
    assign wire3000 = {4'd7, 4'd5};
    assign wire3001 = {4'd7, 4'd5};
    assign wire3002 = {4'd7, 4'd5};
    assign wire3003 = {4'd7, 4'd5};
    assign wire3004 = {4'd7, 4'd5};
    assign wire3005 = {4'd7, 4'd5};
    assign wire3006 = {4'd7, 4'd5};
    assign wire3007 = {4'd7, 4'd5};
    assign wire3008 = {4'd9, 4'd5};
    assign wire3009 = {4'd9, 4'd5};
    assign wire3010 = {4'd9, 4'd5};
    assign wire3011 = {4'd9, 4'd5};
    assign wire3012 = {4'd9, 4'd5};
    assign wire3013 = {4'd11, 4'd7};
    assign wire3014 = {4'd9, 4'd5};
    assign wire3015 = {4'd9, 4'd5};
    assign wire3016 = {4'd10, 4'd6};
    assign wire3017 = {4'd10, 4'd6};
    assign wire3018 = {4'd10, 4'd6};
    assign wire3019 = {4'd10, 4'd6};
    assign wire3020 = {4'd10, 4'd6};
    assign wire3021 = {4'd10, 4'd6};
    assign wire3022 = {4'd10, 4'd6};
    assign wire3023 = {4'd10, 4'd6};
    assign wire3024 = {4'd11, 4'd7};
    assign wire3025 = {4'd11, 4'd7};
    assign wire3026 = {4'd11, 4'd7};
    assign wire3027 = {4'd11, 4'd7};
    assign wire3028 = {4'd11, 4'd7};
    assign wire3029 = {4'd11, 4'd7};
    assign wire3030 = {4'd11, 4'd7};
    assign wire3031 = {4'd11, 4'd7};
    assign wire3032 = {4'd9, 4'd5};
    assign wire3033 = {4'd9, 4'd5};
    assign wire3034 = {4'd9, 4'd5};
    assign wire3035 = {4'd9, 4'd5};
    assign wire3036 = {4'd9, 4'd5};
    assign wire3037 = {4'd9, 4'd5};
    assign wire3038 = {4'd9, 4'd5};
    assign wire3039 = {4'd9, 4'd5};
    assign wire3040 = {4'd11, 4'd5};
    assign wire3041 = {4'd11, 4'd5};
    assign wire3042 = {4'd11, 4'd5};
    assign wire3043 = {4'd11, 4'd5};
    assign wire3044 = {4'd11, 4'd5};
    assign wire3045 = {4'd13, 4'd7};
    assign wire3046 = {4'd11, 4'd5};
    assign wire3047 = {4'd11, 4'd5};
    assign wire3048 = {4'd12, 4'd6};
    assign wire3049 = {4'd12, 4'd6};
    assign wire3050 = {4'd12, 4'd6};
    assign wire3051 = {4'd12, 4'd6};
    assign wire3052 = {4'd12, 4'd6};
    assign wire3053 = {4'd12, 4'd6};
    assign wire3054 = {4'd12, 4'd6};
    assign wire3055 = {4'd12, 4'd6};
    assign wire3056 = {4'd13, 4'd7};
    assign wire3057 = {4'd13, 4'd7};
    assign wire3058 = {4'd13, 4'd7};
    assign wire3059 = {4'd13, 4'd7};
    assign wire3060 = {4'd13, 4'd7};
    assign wire3061 = {4'd13, 4'd7};
    assign wire3062 = {4'd13, 4'd7};
    assign wire3063 = {4'd13, 4'd7};
    assign wire3064 = {4'd11, 4'd5};
    assign wire3065 = {4'd11, 4'd5};
    assign wire3066 = {4'd11, 4'd5};
    assign wire3067 = {4'd11, 4'd5};
    assign wire3068 = {4'd11, 4'd5};
    assign wire3069 = {4'd11, 4'd5};
    assign wire3070 = {4'd11, 4'd5};
    assign wire3071 = {4'd11, 4'd5};
    assign wire3072 = {4'd4, 4'd3};
    assign wire3073 = {4'd4, 4'd3};
    assign wire3074 = {4'd4, 4'd3};
    assign wire3075 = {4'd4, 4'd3};
    assign wire3076 = {4'd4, 4'd3};
    assign wire3077 = {4'd4, 4'd3};
    assign wire3078 = {4'd4, 4'd3};
    assign wire3079 = {4'd4, 4'd3};
    assign wire3080 = {4'd4, 4'd3};
    assign wire3081 = {4'd4, 4'd3};
    assign wire3082 = {4'd4, 4'd3};
    assign wire3083 = {4'd4, 4'd3};
    assign wire3084 = {4'd4, 4'd3};
    assign wire3085 = {4'd4, 4'd3};
    assign wire3086 = {4'd4, 4'd3};
    assign wire3087 = {4'd4, 4'd3};
    assign wire3088 = {4'd4, 4'd3};
    assign wire3089 = {4'd4, 4'd3};
    assign wire3090 = {4'd4, 4'd3};
    assign wire3091 = {4'd4, 4'd3};
    assign wire3092 = {4'd4, 4'd3};
    assign wire3093 = {4'd4, 4'd3};
    assign wire3094 = {4'd4, 4'd3};
    assign wire3095 = {4'd4, 4'd3};
    assign wire3096 = {4'd4, 4'd3};
    assign wire3097 = {4'd4, 4'd3};
    assign wire3098 = {4'd4, 4'd3};
    assign wire3099 = {4'd4, 4'd3};
    assign wire3100 = {4'd4, 4'd3};
    assign wire3101 = {4'd4, 4'd3};
    assign wire3102 = {4'd4, 4'd3};
    assign wire3103 = {4'd4, 4'd3};
    assign wire3104 = {4'd5, 4'd3};
    assign wire3105 = {4'd5, 4'd3};
    assign wire3106 = {4'd5, 4'd3};
    assign wire3107 = {4'd5, 4'd3};
    assign wire3108 = {4'd5, 4'd3};
    assign wire3109 = {4'd5, 4'd3};
    assign wire3110 = {4'd5, 4'd3};
    assign wire3111 = {4'd5, 4'd3};
    assign wire3112 = {4'd5, 4'd3};
    assign wire3113 = {4'd5, 4'd3};
    assign wire3114 = {4'd5, 4'd3};
    assign wire3115 = {4'd5, 4'd3};
    assign wire3116 = {4'd5, 4'd3};
    assign wire3117 = {4'd5, 4'd3};
    assign wire3118 = {4'd5, 4'd3};
    assign wire3119 = {4'd5, 4'd3};
    assign wire3120 = {4'd5, 4'd3};
    assign wire3121 = {4'd5, 4'd3};
    assign wire3122 = {4'd5, 4'd3};
    assign wire3123 = {4'd5, 4'd3};
    assign wire3124 = {4'd5, 4'd3};
    assign wire3125 = {4'd5, 4'd3};
    assign wire3126 = {4'd5, 4'd3};
    assign wire3127 = {4'd5, 4'd3};
    assign wire3128 = {4'd5, 4'd3};
    assign wire3129 = {4'd5, 4'd3};
    assign wire3130 = {4'd5, 4'd3};
    assign wire3131 = {4'd5, 4'd3};
    assign wire3132 = {4'd5, 4'd3};
    assign wire3133 = {4'd5, 4'd3};
    assign wire3134 = {4'd5, 4'd3};
    assign wire3135 = {4'd5, 4'd3};
    assign wire3136 = {4'd7, 4'd3};
    assign wire3137 = {4'd7, 4'd3};
    assign wire3138 = {4'd7, 4'd3};
    assign wire3139 = {4'd7, 4'd3};
    assign wire3140 = {4'd7, 4'd3};
    assign wire3141 = {4'd7, 4'd3};
    assign wire3142 = {4'd7, 4'd3};
    assign wire3143 = {4'd7, 4'd3};
    assign wire3144 = {4'd7, 4'd3};
    assign wire3145 = {4'd7, 4'd3};
    assign wire3146 = {4'd7, 4'd3};
    assign wire3147 = {4'd7, 4'd3};
    assign wire3148 = {4'd7, 4'd3};
    assign wire3149 = {4'd7, 4'd3};
    assign wire3150 = {4'd7, 4'd3};
    assign wire3151 = {4'd7, 4'd3};
    assign wire3152 = {4'd7, 4'd3};
    assign wire3153 = {4'd7, 4'd3};
    assign wire3154 = {4'd7, 4'd3};
    assign wire3155 = {4'd7, 4'd3};
    assign wire3156 = {4'd7, 4'd3};
    assign wire3157 = {4'd7, 4'd3};
    assign wire3158 = {4'd7, 4'd3};
    assign wire3159 = {4'd7, 4'd3};
    assign wire3160 = {4'd7, 4'd3};
    assign wire3161 = {4'd7, 4'd3};
    assign wire3162 = {4'd7, 4'd3};
    assign wire3163 = {4'd7, 4'd3};
    assign wire3164 = {4'd7, 4'd3};
    assign wire3165 = {4'd7, 4'd3};
    assign wire3166 = {4'd7, 4'd3};
    assign wire3167 = {4'd7, 4'd3};
    assign wire3168 = {4'd9, 4'd3};
    assign wire3169 = {4'd9, 4'd3};
    assign wire3170 = {4'd9, 4'd3};
    assign wire3171 = {4'd9, 4'd3};
    assign wire3172 = {4'd9, 4'd3};
    assign wire3173 = {4'd9, 4'd3};
    assign wire3174 = {4'd9, 4'd3};
    assign wire3175 = {4'd9, 4'd3};
    assign wire3176 = {4'd9, 4'd3};
    assign wire3177 = {4'd9, 4'd3};
    assign wire3178 = {4'd9, 4'd3};
    assign wire3179 = {4'd9, 4'd3};
    assign wire3180 = {4'd9, 4'd3};
    assign wire3181 = {4'd9, 4'd3};
    assign wire3182 = {4'd9, 4'd3};
    assign wire3183 = {4'd9, 4'd3};
    assign wire3184 = {4'd9, 4'd3};
    assign wire3185 = {4'd9, 4'd3};
    assign wire3186 = {4'd9, 4'd3};
    assign wire3187 = {4'd9, 4'd3};
    assign wire3188 = {4'd9, 4'd3};
    assign wire3189 = {4'd9, 4'd3};
    assign wire3190 = {4'd9, 4'd3};
    assign wire3191 = {4'd9, 4'd3};
    assign wire3192 = {4'd9, 4'd3};
    assign wire3193 = {4'd9, 4'd3};
    assign wire3194 = {4'd9, 4'd3};
    assign wire3195 = {4'd9, 4'd3};
    assign wire3196 = {4'd9, 4'd3};
    assign wire3197 = {4'd9, 4'd3};
    assign wire3198 = {4'd9, 4'd3};
    assign wire3199 = {4'd9, 4'd3};
    assign wire3200 = {4'd5, 4'd4};
    assign wire3201 = {4'd5, 4'd4};
    assign wire3202 = {4'd5, 4'd4};
    assign wire3203 = {4'd5, 4'd4};
    assign wire3204 = {4'd6, 4'd5};
    assign wire3205 = {4'd9, 4'd8};
    assign wire3206 = {4'd5, 4'd4};
    assign wire3207 = {4'd5, 4'd4};
    assign wire3208 = {4'd6, 4'd5};
    assign wire3209 = {4'd6, 4'd5};
    assign wire3210 = {4'd6, 4'd5};
    assign wire3211 = {4'd6, 4'd5};
    assign wire3212 = {4'd7, 4'd6};
    assign wire3213 = {4'd6, 4'd5};
    assign wire3214 = {4'd6, 4'd5};
    assign wire3215 = {4'd6, 4'd5};
    assign wire3216 = {4'd9, 4'd8};
    assign wire3217 = {4'd9, 4'd8};
    assign wire3218 = {4'd9, 4'd8};
    assign wire3219 = {4'd9, 4'd8};
    assign wire3220 = {4'd10, 4'd9};
    assign wire3221 = {4'd9, 4'd8};
    assign wire3222 = {4'd9, 4'd8};
    assign wire3223 = {4'd9, 4'd8};
    assign wire3224 = {4'd5, 4'd4};
    assign wire3225 = {4'd5, 4'd4};
    assign wire3226 = {4'd5, 4'd4};
    assign wire3227 = {4'd5, 4'd4};
    assign wire3228 = {4'd5, 4'd4};
    assign wire3229 = {4'd5, 4'd4};
    assign wire3230 = {4'd5, 4'd4};
    assign wire3231 = {4'd5, 4'd4};
    assign wire3232 = {4'd6, 4'd4};
    assign wire3233 = {4'd6, 4'd4};
    assign wire3234 = {4'd6, 4'd4};
    assign wire3235 = {4'd6, 4'd4};
    assign wire3236 = {4'd7, 4'd5};
    assign wire3237 = {4'd10, 4'd8};
    assign wire3238 = {4'd6, 4'd4};
    assign wire3239 = {4'd6, 4'd4};
    assign wire3240 = {4'd7, 4'd5};
    assign wire3241 = {4'd7, 4'd5};
    assign wire3242 = {4'd7, 4'd5};
    assign wire3243 = {4'd7, 4'd5};
    assign wire3244 = {4'd8, 4'd6};
    assign wire3245 = {4'd7, 4'd5};
    assign wire3246 = {4'd7, 4'd5};
    assign wire3247 = {4'd7, 4'd5};
    assign wire3248 = {4'd10, 4'd8};
    assign wire3249 = {4'd10, 4'd8};
    assign wire3250 = {4'd10, 4'd8};
    assign wire3251 = {4'd10, 4'd8};
    assign wire3252 = {4'd11, 4'd9};
    assign wire3253 = {4'd10, 4'd8};
    assign wire3254 = {4'd10, 4'd8};
    assign wire3255 = {4'd10, 4'd8};
    assign wire3256 = {4'd6, 4'd4};
    assign wire3257 = {4'd6, 4'd4};
    assign wire3258 = {4'd6, 4'd4};
    assign wire3259 = {4'd6, 4'd4};
    assign wire3260 = {4'd6, 4'd4};
    assign wire3261 = {4'd6, 4'd4};
    assign wire3262 = {4'd6, 4'd4};
    assign wire3263 = {4'd6, 4'd4};
    assign wire3264 = {4'd8, 4'd4};
    assign wire3265 = {4'd8, 4'd4};
    assign wire3266 = {4'd8, 4'd4};
    assign wire3267 = {4'd8, 4'd4};
    assign wire3268 = {4'd9, 4'd5};
    assign wire3269 = {4'd12, 4'd8};
    assign wire3270 = {4'd8, 4'd4};
    assign wire3271 = {4'd8, 4'd4};
    assign wire3272 = {4'd9, 4'd5};
    assign wire3273 = {4'd9, 4'd5};
    assign wire3274 = {4'd9, 4'd5};
    assign wire3275 = {4'd9, 4'd5};
    assign wire3276 = {4'd10, 4'd6};
    assign wire3277 = {4'd9, 4'd5};
    assign wire3278 = {4'd9, 4'd5};
    assign wire3279 = {4'd9, 4'd5};
    assign wire3280 = {4'd12, 4'd8};
    assign wire3281 = {4'd12, 4'd8};
    assign wire3282 = {4'd12, 4'd8};
    assign wire3283 = {4'd12, 4'd8};
    assign wire3284 = {4'd13, 4'd9};
    assign wire3285 = {4'd12, 4'd8};
    assign wire3286 = {4'd12, 4'd8};
    assign wire3287 = {4'd12, 4'd8};
    assign wire3288 = {4'd8, 4'd4};
    assign wire3289 = {4'd8, 4'd4};
    assign wire3290 = {4'd8, 4'd4};
    assign wire3291 = {4'd8, 4'd4};
    assign wire3292 = {4'd8, 4'd4};
    assign wire3293 = {4'd8, 4'd4};
    assign wire3294 = {4'd8, 4'd4};
    assign wire3295 = {4'd8, 4'd4};
    assign wire3296 = {4'd10, 4'd4};
    assign wire3297 = {4'd10, 4'd4};
    assign wire3298 = {4'd10, 4'd4};
    assign wire3299 = {4'd10, 4'd4};
    assign wire3300 = {4'd11, 4'd5};
    assign wire3301 = {4'd14, 4'd8};
    assign wire3302 = {4'd10, 4'd4};
    assign wire3303 = {4'd10, 4'd4};
    assign wire3304 = {4'd11, 4'd5};
    assign wire3305 = {4'd11, 4'd5};
    assign wire3306 = {4'd11, 4'd5};
    assign wire3307 = {4'd11, 4'd5};
    assign wire3308 = {4'd12, 4'd6};
    assign wire3309 = {4'd11, 4'd5};
    assign wire3310 = {4'd11, 4'd5};
    assign wire3311 = {4'd11, 4'd5};
    assign wire3312 = {4'd14, 4'd8};
    assign wire3313 = {4'd14, 4'd8};
    assign wire3314 = {4'd14, 4'd8};
    assign wire3315 = {4'd14, 4'd8};
    assign wire3316 = {4'd15, 4'd9};
    assign wire3317 = {4'd14, 4'd8};
    assign wire3318 = {4'd14, 4'd8};
    assign wire3319 = {4'd14, 4'd8};
    assign wire3320 = {4'd10, 4'd4};
    assign wire3321 = {4'd10, 4'd4};
    assign wire3322 = {4'd10, 4'd4};
    assign wire3323 = {4'd10, 4'd4};
    assign wire3324 = {4'd10, 4'd4};
    assign wire3325 = {4'd10, 4'd4};
    assign wire3326 = {4'd10, 4'd4};
    assign wire3327 = {4'd10, 4'd4};
    assign wire3328 = {4'd5, 4'd4};
    assign wire3329 = {4'd5, 4'd4};
    assign wire3330 = {4'd5, 4'd4};
    assign wire3331 = {4'd5, 4'd4};
    assign wire3332 = {4'd5, 4'd4};
    assign wire3333 = {4'd5, 4'd4};
    assign wire3334 = {4'd5, 4'd4};
    assign wire3335 = {4'd5, 4'd4};
    assign wire3336 = {4'd5, 4'd4};
    assign wire3337 = {4'd5, 4'd4};
    assign wire3338 = {4'd5, 4'd4};
    assign wire3339 = {4'd5, 4'd4};
    assign wire3340 = {4'd5, 4'd4};
    assign wire3341 = {4'd5, 4'd4};
    assign wire3342 = {4'd5, 4'd4};
    assign wire3343 = {4'd5, 4'd4};
    assign wire3344 = {4'd5, 4'd4};
    assign wire3345 = {4'd5, 4'd4};
    assign wire3346 = {4'd5, 4'd4};
    assign wire3347 = {4'd5, 4'd4};
    assign wire3348 = {4'd5, 4'd4};
    assign wire3349 = {4'd5, 4'd4};
    assign wire3350 = {4'd5, 4'd4};
    assign wire3351 = {4'd5, 4'd4};
    assign wire3352 = {4'd5, 4'd4};
    assign wire3353 = {4'd5, 4'd4};
    assign wire3354 = {4'd5, 4'd4};
    assign wire3355 = {4'd5, 4'd4};
    assign wire3356 = {4'd5, 4'd4};
    assign wire3357 = {4'd5, 4'd4};
    assign wire3358 = {4'd5, 4'd4};
    assign wire3359 = {4'd5, 4'd4};
    assign wire3360 = {4'd6, 4'd4};
    assign wire3361 = {4'd6, 4'd4};
    assign wire3362 = {4'd6, 4'd4};
    assign wire3363 = {4'd6, 4'd4};
    assign wire3364 = {4'd6, 4'd4};
    assign wire3365 = {4'd6, 4'd4};
    assign wire3366 = {4'd6, 4'd4};
    assign wire3367 = {4'd6, 4'd4};
    assign wire3368 = {4'd6, 4'd4};
    assign wire3369 = {4'd6, 4'd4};
    assign wire3370 = {4'd6, 4'd4};
    assign wire3371 = {4'd6, 4'd4};
    assign wire3372 = {4'd6, 4'd4};
    assign wire3373 = {4'd6, 4'd4};
    assign wire3374 = {4'd6, 4'd4};
    assign wire3375 = {4'd6, 4'd4};
    assign wire3376 = {4'd6, 4'd4};
    assign wire3377 = {4'd6, 4'd4};
    assign wire3378 = {4'd6, 4'd4};
    assign wire3379 = {4'd6, 4'd4};
    assign wire3380 = {4'd6, 4'd4};
    assign wire3381 = {4'd6, 4'd4};
    assign wire3382 = {4'd6, 4'd4};
    assign wire3383 = {4'd6, 4'd4};
    assign wire3384 = {4'd6, 4'd4};
    assign wire3385 = {4'd6, 4'd4};
    assign wire3386 = {4'd6, 4'd4};
    assign wire3387 = {4'd6, 4'd4};
    assign wire3388 = {4'd6, 4'd4};
    assign wire3389 = {4'd6, 4'd4};
    assign wire3390 = {4'd6, 4'd4};
    assign wire3391 = {4'd6, 4'd4};
    assign wire3392 = {4'd8, 4'd4};
    assign wire3393 = {4'd8, 4'd4};
    assign wire3394 = {4'd8, 4'd4};
    assign wire3395 = {4'd8, 4'd4};
    assign wire3396 = {4'd8, 4'd4};
    assign wire3397 = {4'd8, 4'd4};
    assign wire3398 = {4'd8, 4'd4};
    assign wire3399 = {4'd8, 4'd4};
    assign wire3400 = {4'd8, 4'd4};
    assign wire3401 = {4'd8, 4'd4};
    assign wire3402 = {4'd8, 4'd4};
    assign wire3403 = {4'd8, 4'd4};
    assign wire3404 = {4'd8, 4'd4};
    assign wire3405 = {4'd8, 4'd4};
    assign wire3406 = {4'd8, 4'd4};
    assign wire3407 = {4'd8, 4'd4};
    assign wire3408 = {4'd8, 4'd4};
    assign wire3409 = {4'd8, 4'd4};
    assign wire3410 = {4'd8, 4'd4};
    assign wire3411 = {4'd8, 4'd4};
    assign wire3412 = {4'd8, 4'd4};
    assign wire3413 = {4'd8, 4'd4};
    assign wire3414 = {4'd8, 4'd4};
    assign wire3415 = {4'd8, 4'd4};
    assign wire3416 = {4'd8, 4'd4};
    assign wire3417 = {4'd8, 4'd4};
    assign wire3418 = {4'd8, 4'd4};
    assign wire3419 = {4'd8, 4'd4};
    assign wire3420 = {4'd8, 4'd4};
    assign wire3421 = {4'd8, 4'd4};
    assign wire3422 = {4'd8, 4'd4};
    assign wire3423 = {4'd8, 4'd4};
    assign wire3424 = {4'd10, 4'd4};
    assign wire3425 = {4'd10, 4'd4};
    assign wire3426 = {4'd10, 4'd4};
    assign wire3427 = {4'd10, 4'd4};
    assign wire3428 = {4'd10, 4'd4};
    assign wire3429 = {4'd10, 4'd4};
    assign wire3430 = {4'd10, 4'd4};
    assign wire3431 = {4'd10, 4'd4};
    assign wire3432 = {4'd10, 4'd4};
    assign wire3433 = {4'd10, 4'd4};
    assign wire3434 = {4'd10, 4'd4};
    assign wire3435 = {4'd10, 4'd4};
    assign wire3436 = {4'd10, 4'd4};
    assign wire3437 = {4'd10, 4'd4};
    assign wire3438 = {4'd10, 4'd4};
    assign wire3439 = {4'd10, 4'd4};
    assign wire3440 = {4'd10, 4'd4};
    assign wire3441 = {4'd10, 4'd4};
    assign wire3442 = {4'd10, 4'd4};
    assign wire3443 = {4'd10, 4'd4};
    assign wire3444 = {4'd10, 4'd4};
    assign wire3445 = {4'd10, 4'd4};
    assign wire3446 = {4'd10, 4'd4};
    assign wire3447 = {4'd10, 4'd4};
    assign wire3448 = {4'd10, 4'd4};
    assign wire3449 = {4'd10, 4'd4};
    assign wire3450 = {4'd10, 4'd4};
    assign wire3451 = {4'd10, 4'd4};
    assign wire3452 = {4'd10, 4'd4};
    assign wire3453 = {4'd10, 4'd4};
    assign wire3454 = {4'd10, 4'd4};
    assign wire3455 = {4'd10, 4'd4};
    assign wire3456 = {4'd6, 4'd5};
    assign wire3457 = {4'd6, 4'd5};
    assign wire3458 = {4'd6, 4'd5};
    assign wire3459 = {4'd6, 4'd5};
    assign wire3460 = {4'd7, 4'd6};
    assign wire3461 = {4'd10, 4'd9};
    assign wire3462 = {4'd6, 4'd5};
    assign wire3463 = {4'd6, 4'd5};
    assign wire3464 = {4'd7, 4'd6};
    assign wire3465 = {4'd7, 4'd6};
    assign wire3466 = {4'd7, 4'd6};
    assign wire3467 = {4'd7, 4'd6};
    assign wire3468 = {4'd8, 4'd7};
    assign wire3469 = {4'd7, 4'd6};
    assign wire3470 = {4'd7, 4'd6};
    assign wire3471 = {4'd7, 4'd6};
    assign wire3472 = {4'd10, 4'd9};
    assign wire3473 = {4'd10, 4'd9};
    assign wire3474 = {4'd10, 4'd9};
    assign wire3475 = {4'd10, 4'd9};
    assign wire3476 = {4'd11, 4'd10};
    assign wire3477 = {4'd10, 4'd9};
    assign wire3478 = {4'd10, 4'd9};
    assign wire3479 = {4'd10, 4'd9};
    assign wire3480 = {4'd6, 4'd5};
    assign wire3481 = {4'd6, 4'd5};
    assign wire3482 = {4'd6, 4'd5};
    assign wire3483 = {4'd6, 4'd5};
    assign wire3484 = {4'd6, 4'd5};
    assign wire3485 = {4'd6, 4'd5};
    assign wire3486 = {4'd6, 4'd5};
    assign wire3487 = {4'd6, 4'd5};
    assign wire3488 = {4'd7, 4'd5};
    assign wire3489 = {4'd7, 4'd5};
    assign wire3490 = {4'd7, 4'd5};
    assign wire3491 = {4'd7, 4'd5};
    assign wire3492 = {4'd8, 4'd6};
    assign wire3493 = {4'd11, 4'd9};
    assign wire3494 = {4'd7, 4'd5};
    assign wire3495 = {4'd7, 4'd5};
    assign wire3496 = {4'd8, 4'd6};
    assign wire3497 = {4'd8, 4'd6};
    assign wire3498 = {4'd8, 4'd6};
    assign wire3499 = {4'd8, 4'd6};
    assign wire3500 = {4'd9, 4'd7};
    assign wire3501 = {4'd8, 4'd6};
    assign wire3502 = {4'd8, 4'd6};
    assign wire3503 = {4'd8, 4'd6};
    assign wire3504 = {4'd11, 4'd9};
    assign wire3505 = {4'd11, 4'd9};
    assign wire3506 = {4'd11, 4'd9};
    assign wire3507 = {4'd11, 4'd9};
    assign wire3508 = {4'd12, 4'd10};
    assign wire3509 = {4'd11, 4'd9};
    assign wire3510 = {4'd11, 4'd9};
    assign wire3511 = {4'd11, 4'd9};
    assign wire3512 = {4'd7, 4'd5};
    assign wire3513 = {4'd7, 4'd5};
    assign wire3514 = {4'd7, 4'd5};
    assign wire3515 = {4'd7, 4'd5};
    assign wire3516 = {4'd7, 4'd5};
    assign wire3517 = {4'd7, 4'd5};
    assign wire3518 = {4'd7, 4'd5};
    assign wire3519 = {4'd7, 4'd5};
    assign wire3520 = {4'd9, 4'd5};
    assign wire3521 = {4'd9, 4'd5};
    assign wire3522 = {4'd9, 4'd5};
    assign wire3523 = {4'd9, 4'd5};
    assign wire3524 = {4'd10, 4'd6};
    assign wire3525 = {4'd13, 4'd9};
    assign wire3526 = {4'd9, 4'd5};
    assign wire3527 = {4'd9, 4'd5};
    assign wire3528 = {4'd10, 4'd6};
    assign wire3529 = {4'd10, 4'd6};
    assign wire3530 = {4'd10, 4'd6};
    assign wire3531 = {4'd10, 4'd6};
    assign wire3532 = {4'd11, 4'd7};
    assign wire3533 = {4'd10, 4'd6};
    assign wire3534 = {4'd10, 4'd6};
    assign wire3535 = {4'd10, 4'd6};
    assign wire3536 = {4'd13, 4'd9};
    assign wire3537 = {4'd13, 4'd9};
    assign wire3538 = {4'd13, 4'd9};
    assign wire3539 = {4'd13, 4'd9};
    assign wire3540 = {4'd14, 4'd10};
    assign wire3541 = {4'd13, 4'd9};
    assign wire3542 = {4'd13, 4'd9};
    assign wire3543 = {4'd13, 4'd9};
    assign wire3544 = {4'd9, 4'd5};
    assign wire3545 = {4'd9, 4'd5};
    assign wire3546 = {4'd9, 4'd5};
    assign wire3547 = {4'd9, 4'd5};
    assign wire3548 = {4'd9, 4'd5};
    assign wire3549 = {4'd9, 4'd5};
    assign wire3550 = {4'd9, 4'd5};
    assign wire3551 = {4'd9, 4'd5};
    assign wire3552 = {4'd11, 4'd5};
    assign wire3553 = {4'd11, 4'd5};
    assign wire3554 = {4'd11, 4'd5};
    assign wire3555 = {4'd11, 4'd5};
    assign wire3556 = {4'd12, 4'd6};
    assign wire3557 = {4'd15, 4'd9};
    assign wire3558 = {4'd11, 4'd5};
    assign wire3559 = {4'd11, 4'd5};
    assign wire3560 = {4'd12, 4'd6};
    assign wire3561 = {4'd12, 4'd6};
    assign wire3562 = {4'd12, 4'd6};
    assign wire3563 = {4'd12, 4'd6};
    assign wire3564 = {4'd13, 4'd7};
    assign wire3565 = {4'd12, 4'd6};
    assign wire3566 = {4'd12, 4'd6};
    assign wire3567 = {4'd12, 4'd6};
    assign wire3568 = {4'd15, 4'd9};
    assign wire3569 = {4'd15, 4'd9};
    assign wire3570 = {4'd15, 4'd9};
    assign wire3571 = {4'd15, 4'd9};
    assign wire3572 = {4'd16, 4'd10};
    assign wire3573 = {4'd15, 4'd9};
    assign wire3574 = {4'd15, 4'd9};
    assign wire3575 = {4'd15, 4'd9};
    assign wire3576 = {4'd11, 4'd5};
    assign wire3577 = {4'd11, 4'd5};
    assign wire3578 = {4'd11, 4'd5};
    assign wire3579 = {4'd11, 4'd5};
    assign wire3580 = {4'd11, 4'd5};
    assign wire3581 = {4'd11, 4'd5};
    assign wire3582 = {4'd11, 4'd5};
    assign wire3583 = {4'd11, 4'd5};
    assign wire3584 = {4'd5, 4'd4};
    assign wire3585 = {4'd5, 4'd4};
    assign wire3586 = {4'd5, 4'd4};
    assign wire3587 = {4'd5, 4'd4};
    assign wire3588 = {4'd5, 4'd4};
    assign wire3589 = {4'd5, 4'd4};
    assign wire3590 = {4'd5, 4'd4};
    assign wire3591 = {4'd5, 4'd4};
    assign wire3592 = {4'd5, 4'd4};
    assign wire3593 = {4'd5, 4'd4};
    assign wire3594 = {4'd5, 4'd4};
    assign wire3595 = {4'd5, 4'd4};
    assign wire3596 = {4'd5, 4'd4};
    assign wire3597 = {4'd5, 4'd4};
    assign wire3598 = {4'd5, 4'd4};
    assign wire3599 = {4'd5, 4'd4};
    assign wire3600 = {4'd5, 4'd4};
    assign wire3601 = {4'd5, 4'd4};
    assign wire3602 = {4'd5, 4'd4};
    assign wire3603 = {4'd5, 4'd4};
    assign wire3604 = {4'd5, 4'd4};
    assign wire3605 = {4'd5, 4'd4};
    assign wire3606 = {4'd5, 4'd4};
    assign wire3607 = {4'd5, 4'd4};
    assign wire3608 = {4'd5, 4'd4};
    assign wire3609 = {4'd5, 4'd4};
    assign wire3610 = {4'd5, 4'd4};
    assign wire3611 = {4'd5, 4'd4};
    assign wire3612 = {4'd5, 4'd4};
    assign wire3613 = {4'd5, 4'd4};
    assign wire3614 = {4'd5, 4'd4};
    assign wire3615 = {4'd5, 4'd4};
    assign wire3616 = {4'd6, 4'd4};
    assign wire3617 = {4'd6, 4'd4};
    assign wire3618 = {4'd6, 4'd4};
    assign wire3619 = {4'd6, 4'd4};
    assign wire3620 = {4'd6, 4'd4};
    assign wire3621 = {4'd6, 4'd4};
    assign wire3622 = {4'd6, 4'd4};
    assign wire3623 = {4'd6, 4'd4};
    assign wire3624 = {4'd6, 4'd4};
    assign wire3625 = {4'd6, 4'd4};
    assign wire3626 = {4'd6, 4'd4};
    assign wire3627 = {4'd6, 4'd4};
    assign wire3628 = {4'd6, 4'd4};
    assign wire3629 = {4'd6, 4'd4};
    assign wire3630 = {4'd6, 4'd4};
    assign wire3631 = {4'd6, 4'd4};
    assign wire3632 = {4'd6, 4'd4};
    assign wire3633 = {4'd6, 4'd4};
    assign wire3634 = {4'd6, 4'd4};
    assign wire3635 = {4'd6, 4'd4};
    assign wire3636 = {4'd6, 4'd4};
    assign wire3637 = {4'd6, 4'd4};
    assign wire3638 = {4'd6, 4'd4};
    assign wire3639 = {4'd6, 4'd4};
    assign wire3640 = {4'd6, 4'd4};
    assign wire3641 = {4'd6, 4'd4};
    assign wire3642 = {4'd6, 4'd4};
    assign wire3643 = {4'd6, 4'd4};
    assign wire3644 = {4'd6, 4'd4};
    assign wire3645 = {4'd6, 4'd4};
    assign wire3646 = {4'd6, 4'd4};
    assign wire3647 = {4'd6, 4'd4};
    assign wire3648 = {4'd8, 4'd4};
    assign wire3649 = {4'd8, 4'd4};
    assign wire3650 = {4'd8, 4'd4};
    assign wire3651 = {4'd8, 4'd4};
    assign wire3652 = {4'd8, 4'd4};
    assign wire3653 = {4'd8, 4'd4};
    assign wire3654 = {4'd8, 4'd4};
    assign wire3655 = {4'd8, 4'd4};
    assign wire3656 = {4'd8, 4'd4};
    assign wire3657 = {4'd8, 4'd4};
    assign wire3658 = {4'd8, 4'd4};
    assign wire3659 = {4'd8, 4'd4};
    assign wire3660 = {4'd8, 4'd4};
    assign wire3661 = {4'd8, 4'd4};
    assign wire3662 = {4'd8, 4'd4};
    assign wire3663 = {4'd8, 4'd4};
    assign wire3664 = {4'd8, 4'd4};
    assign wire3665 = {4'd8, 4'd4};
    assign wire3666 = {4'd8, 4'd4};
    assign wire3667 = {4'd8, 4'd4};
    assign wire3668 = {4'd8, 4'd4};
    assign wire3669 = {4'd8, 4'd4};
    assign wire3670 = {4'd8, 4'd4};
    assign wire3671 = {4'd8, 4'd4};
    assign wire3672 = {4'd8, 4'd4};
    assign wire3673 = {4'd8, 4'd4};
    assign wire3674 = {4'd8, 4'd4};
    assign wire3675 = {4'd8, 4'd4};
    assign wire3676 = {4'd8, 4'd4};
    assign wire3677 = {4'd8, 4'd4};
    assign wire3678 = {4'd8, 4'd4};
    assign wire3679 = {4'd8, 4'd4};
    assign wire3680 = {4'd10, 4'd4};
    assign wire3681 = {4'd10, 4'd4};
    assign wire3682 = {4'd10, 4'd4};
    assign wire3683 = {4'd10, 4'd4};
    assign wire3684 = {4'd10, 4'd4};
    assign wire3685 = {4'd10, 4'd4};
    assign wire3686 = {4'd10, 4'd4};
    assign wire3687 = {4'd10, 4'd4};
    assign wire3688 = {4'd10, 4'd4};
    assign wire3689 = {4'd10, 4'd4};
    assign wire3690 = {4'd10, 4'd4};
    assign wire3691 = {4'd10, 4'd4};
    assign wire3692 = {4'd10, 4'd4};
    assign wire3693 = {4'd10, 4'd4};
    assign wire3694 = {4'd10, 4'd4};
    assign wire3695 = {4'd10, 4'd4};
    assign wire3696 = {4'd10, 4'd4};
    assign wire3697 = {4'd10, 4'd4};
    assign wire3698 = {4'd10, 4'd4};
    assign wire3699 = {4'd10, 4'd4};
    assign wire3700 = {4'd10, 4'd4};
    assign wire3701 = {4'd10, 4'd4};
    assign wire3702 = {4'd10, 4'd4};
    assign wire3703 = {4'd10, 4'd4};
    assign wire3704 = {4'd10, 4'd4};
    assign wire3705 = {4'd10, 4'd4};
    assign wire3706 = {4'd10, 4'd4};
    assign wire3707 = {4'd10, 4'd4};
    assign wire3708 = {4'd10, 4'd4};
    assign wire3709 = {4'd10, 4'd4};
    assign wire3710 = {4'd10, 4'd4};
    assign wire3711 = {4'd10, 4'd4};
    assign wire3712 = {4'd6, 4'd5};
    assign wire3713 = {4'd6, 4'd5};
    assign wire3714 = {4'd6, 4'd5};
    assign wire3715 = {4'd6, 4'd5};
    assign wire3716 = {4'd6, 4'd5};
    assign wire3717 = {4'd8, 4'd7};
    assign wire3718 = {4'd6, 4'd5};
    assign wire3719 = {4'd6, 4'd5};
    assign wire3720 = {4'd7, 4'd6};
    assign wire3721 = {4'd7, 4'd6};
    assign wire3722 = {4'd7, 4'd6};
    assign wire3723 = {4'd7, 4'd6};
    assign wire3724 = {4'd7, 4'd6};
    assign wire3725 = {4'd7, 4'd6};
    assign wire3726 = {4'd7, 4'd6};
    assign wire3727 = {4'd7, 4'd6};
    assign wire3728 = {4'd8, 4'd7};
    assign wire3729 = {4'd8, 4'd7};
    assign wire3730 = {4'd8, 4'd7};
    assign wire3731 = {4'd8, 4'd7};
    assign wire3732 = {4'd8, 4'd7};
    assign wire3733 = {4'd8, 4'd7};
    assign wire3734 = {4'd8, 4'd7};
    assign wire3735 = {4'd8, 4'd7};
    assign wire3736 = {4'd6, 4'd5};
    assign wire3737 = {4'd6, 4'd5};
    assign wire3738 = {4'd6, 4'd5};
    assign wire3739 = {4'd6, 4'd5};
    assign wire3740 = {4'd6, 4'd5};
    assign wire3741 = {4'd6, 4'd5};
    assign wire3742 = {4'd6, 4'd5};
    assign wire3743 = {4'd6, 4'd5};
    assign wire3744 = {4'd7, 4'd5};
    assign wire3745 = {4'd7, 4'd5};
    assign wire3746 = {4'd7, 4'd5};
    assign wire3747 = {4'd7, 4'd5};
    assign wire3748 = {4'd7, 4'd5};
    assign wire3749 = {4'd9, 4'd7};
    assign wire3750 = {4'd7, 4'd5};
    assign wire3751 = {4'd7, 4'd5};
    assign wire3752 = {4'd8, 4'd6};
    assign wire3753 = {4'd8, 4'd6};
    assign wire3754 = {4'd8, 4'd6};
    assign wire3755 = {4'd8, 4'd6};
    assign wire3756 = {4'd8, 4'd6};
    assign wire3757 = {4'd8, 4'd6};
    assign wire3758 = {4'd8, 4'd6};
    assign wire3759 = {4'd8, 4'd6};
    assign wire3760 = {4'd9, 4'd7};
    assign wire3761 = {4'd9, 4'd7};
    assign wire3762 = {4'd9, 4'd7};
    assign wire3763 = {4'd9, 4'd7};
    assign wire3764 = {4'd9, 4'd7};
    assign wire3765 = {4'd9, 4'd7};
    assign wire3766 = {4'd9, 4'd7};
    assign wire3767 = {4'd9, 4'd7};
    assign wire3768 = {4'd7, 4'd5};
    assign wire3769 = {4'd7, 4'd5};
    assign wire3770 = {4'd7, 4'd5};
    assign wire3771 = {4'd7, 4'd5};
    assign wire3772 = {4'd7, 4'd5};
    assign wire3773 = {4'd7, 4'd5};
    assign wire3774 = {4'd7, 4'd5};
    assign wire3775 = {4'd7, 4'd5};
    assign wire3776 = {4'd9, 4'd5};
    assign wire3777 = {4'd9, 4'd5};
    assign wire3778 = {4'd9, 4'd5};
    assign wire3779 = {4'd9, 4'd5};
    assign wire3780 = {4'd9, 4'd5};
    assign wire3781 = {4'd11, 4'd7};
    assign wire3782 = {4'd9, 4'd5};
    assign wire3783 = {4'd9, 4'd5};
    assign wire3784 = {4'd10, 4'd6};
    assign wire3785 = {4'd10, 4'd6};
    assign wire3786 = {4'd10, 4'd6};
    assign wire3787 = {4'd10, 4'd6};
    assign wire3788 = {4'd10, 4'd6};
    assign wire3789 = {4'd10, 4'd6};
    assign wire3790 = {4'd10, 4'd6};
    assign wire3791 = {4'd10, 4'd6};
    assign wire3792 = {4'd11, 4'd7};
    assign wire3793 = {4'd11, 4'd7};
    assign wire3794 = {4'd11, 4'd7};
    assign wire3795 = {4'd11, 4'd7};
    assign wire3796 = {4'd11, 4'd7};
    assign wire3797 = {4'd11, 4'd7};
    assign wire3798 = {4'd11, 4'd7};
    assign wire3799 = {4'd11, 4'd7};
    assign wire3800 = {4'd9, 4'd5};
    assign wire3801 = {4'd9, 4'd5};
    assign wire3802 = {4'd9, 4'd5};
    assign wire3803 = {4'd9, 4'd5};
    assign wire3804 = {4'd9, 4'd5};
    assign wire3805 = {4'd9, 4'd5};
    assign wire3806 = {4'd9, 4'd5};
    assign wire3807 = {4'd9, 4'd5};
    assign wire3808 = {4'd11, 4'd5};
    assign wire3809 = {4'd11, 4'd5};
    assign wire3810 = {4'd11, 4'd5};
    assign wire3811 = {4'd11, 4'd5};
    assign wire3812 = {4'd11, 4'd5};
    assign wire3813 = {4'd13, 4'd7};
    assign wire3814 = {4'd11, 4'd5};
    assign wire3815 = {4'd11, 4'd5};
    assign wire3816 = {4'd12, 4'd6};
    assign wire3817 = {4'd12, 4'd6};
    assign wire3818 = {4'd12, 4'd6};
    assign wire3819 = {4'd12, 4'd6};
    assign wire3820 = {4'd12, 4'd6};
    assign wire3821 = {4'd12, 4'd6};
    assign wire3822 = {4'd12, 4'd6};
    assign wire3823 = {4'd12, 4'd6};
    assign wire3824 = {4'd13, 4'd7};
    assign wire3825 = {4'd13, 4'd7};
    assign wire3826 = {4'd13, 4'd7};
    assign wire3827 = {4'd13, 4'd7};
    assign wire3828 = {4'd13, 4'd7};
    assign wire3829 = {4'd13, 4'd7};
    assign wire3830 = {4'd13, 4'd7};
    assign wire3831 = {4'd13, 4'd7};
    assign wire3832 = {4'd11, 4'd5};
    assign wire3833 = {4'd11, 4'd5};
    assign wire3834 = {4'd11, 4'd5};
    assign wire3835 = {4'd11, 4'd5};
    assign wire3836 = {4'd11, 4'd5};
    assign wire3837 = {4'd11, 4'd5};
    assign wire3838 = {4'd11, 4'd5};
    assign wire3839 = {4'd11, 4'd5};
    assign wire3840 = {4'd6, 4'd5};
    assign wire3841 = {4'd6, 4'd5};
    assign wire3842 = {4'd6, 4'd5};
    assign wire3843 = {4'd6, 4'd5};
    assign wire3844 = {4'd6, 4'd5};
    assign wire3845 = {4'd6, 4'd5};
    assign wire3846 = {4'd6, 4'd5};
    assign wire3847 = {4'd6, 4'd5};
    assign wire3848 = {4'd6, 4'd5};
    assign wire3849 = {4'd6, 4'd5};
    assign wire3850 = {4'd6, 4'd5};
    assign wire3851 = {4'd6, 4'd5};
    assign wire3852 = {4'd6, 4'd5};
    assign wire3853 = {4'd6, 4'd5};
    assign wire3854 = {4'd6, 4'd5};
    assign wire3855 = {4'd6, 4'd5};
    assign wire3856 = {4'd6, 4'd5};
    assign wire3857 = {4'd6, 4'd5};
    assign wire3858 = {4'd6, 4'd5};
    assign wire3859 = {4'd6, 4'd5};
    assign wire3860 = {4'd6, 4'd5};
    assign wire3861 = {4'd6, 4'd5};
    assign wire3862 = {4'd6, 4'd5};
    assign wire3863 = {4'd6, 4'd5};
    assign wire3864 = {4'd6, 4'd5};
    assign wire3865 = {4'd6, 4'd5};
    assign wire3866 = {4'd6, 4'd5};
    assign wire3867 = {4'd6, 4'd5};
    assign wire3868 = {4'd6, 4'd5};
    assign wire3869 = {4'd6, 4'd5};
    assign wire3870 = {4'd6, 4'd5};
    assign wire3871 = {4'd6, 4'd5};
    assign wire3872 = {4'd7, 4'd5};
    assign wire3873 = {4'd7, 4'd5};
    assign wire3874 = {4'd7, 4'd5};
    assign wire3875 = {4'd7, 4'd5};
    assign wire3876 = {4'd7, 4'd5};
    assign wire3877 = {4'd7, 4'd5};
    assign wire3878 = {4'd7, 4'd5};
    assign wire3879 = {4'd7, 4'd5};
    assign wire3880 = {4'd7, 4'd5};
    assign wire3881 = {4'd7, 4'd5};
    assign wire3882 = {4'd7, 4'd5};
    assign wire3883 = {4'd7, 4'd5};
    assign wire3884 = {4'd7, 4'd5};
    assign wire3885 = {4'd7, 4'd5};
    assign wire3886 = {4'd7, 4'd5};
    assign wire3887 = {4'd7, 4'd5};
    assign wire3888 = {4'd7, 4'd5};
    assign wire3889 = {4'd7, 4'd5};
    assign wire3890 = {4'd7, 4'd5};
    assign wire3891 = {4'd7, 4'd5};
    assign wire3892 = {4'd7, 4'd5};
    assign wire3893 = {4'd7, 4'd5};
    assign wire3894 = {4'd7, 4'd5};
    assign wire3895 = {4'd7, 4'd5};
    assign wire3896 = {4'd7, 4'd5};
    assign wire3897 = {4'd7, 4'd5};
    assign wire3898 = {4'd7, 4'd5};
    assign wire3899 = {4'd7, 4'd5};
    assign wire3900 = {4'd7, 4'd5};
    assign wire3901 = {4'd7, 4'd5};
    assign wire3902 = {4'd7, 4'd5};
    assign wire3903 = {4'd7, 4'd5};
    assign wire3904 = {4'd9, 4'd5};
    assign wire3905 = {4'd9, 4'd5};
    assign wire3906 = {4'd9, 4'd5};
    assign wire3907 = {4'd9, 4'd5};
    assign wire3908 = {4'd9, 4'd5};
    assign wire3909 = {4'd9, 4'd5};
    assign wire3910 = {4'd9, 4'd5};
    assign wire3911 = {4'd9, 4'd5};
    assign wire3912 = {4'd9, 4'd5};
    assign wire3913 = {4'd9, 4'd5};
    assign wire3914 = {4'd9, 4'd5};
    assign wire3915 = {4'd9, 4'd5};
    assign wire3916 = {4'd9, 4'd5};
    assign wire3917 = {4'd9, 4'd5};
    assign wire3918 = {4'd9, 4'd5};
    assign wire3919 = {4'd9, 4'd5};
    assign wire3920 = {4'd9, 4'd5};
    assign wire3921 = {4'd9, 4'd5};
    assign wire3922 = {4'd9, 4'd5};
    assign wire3923 = {4'd9, 4'd5};
    assign wire3924 = {4'd9, 4'd5};
    assign wire3925 = {4'd9, 4'd5};
    assign wire3926 = {4'd9, 4'd5};
    assign wire3927 = {4'd9, 4'd5};
    assign wire3928 = {4'd9, 4'd5};
    assign wire3929 = {4'd9, 4'd5};
    assign wire3930 = {4'd9, 4'd5};
    assign wire3931 = {4'd9, 4'd5};
    assign wire3932 = {4'd9, 4'd5};
    assign wire3933 = {4'd9, 4'd5};
    assign wire3934 = {4'd9, 4'd5};
    assign wire3935 = {4'd9, 4'd5};
    assign wire3936 = {4'd11, 4'd5};
    assign wire3937 = {4'd11, 4'd5};
    assign wire3938 = {4'd11, 4'd5};
    assign wire3939 = {4'd11, 4'd5};
    assign wire3940 = {4'd11, 4'd5};
    assign wire3941 = {4'd11, 4'd5};
    assign wire3942 = {4'd11, 4'd5};
    assign wire3943 = {4'd11, 4'd5};
    assign wire3944 = {4'd11, 4'd5};
    assign wire3945 = {4'd11, 4'd5};
    assign wire3946 = {4'd11, 4'd5};
    assign wire3947 = {4'd11, 4'd5};
    assign wire3948 = {4'd11, 4'd5};
    assign wire3949 = {4'd11, 4'd5};
    assign wire3950 = {4'd11, 4'd5};
    assign wire3951 = {4'd11, 4'd5};
    assign wire3952 = {4'd11, 4'd5};
    assign wire3953 = {4'd11, 4'd5};
    assign wire3954 = {4'd11, 4'd5};
    assign wire3955 = {4'd11, 4'd5};
    assign wire3956 = {4'd11, 4'd5};
    assign wire3957 = {4'd11, 4'd5};
    assign wire3958 = {4'd11, 4'd5};
    assign wire3959 = {4'd11, 4'd5};
    assign wire3960 = {4'd11, 4'd5};
    assign wire3961 = {4'd11, 4'd5};
    assign wire3962 = {4'd11, 4'd5};
    assign wire3963 = {4'd11, 4'd5};
    assign wire3964 = {4'd11, 4'd5};
    assign wire3965 = {4'd11, 4'd5};
    assign wire3966 = {4'd11, 4'd5};
    assign wire3967 = {4'd11, 4'd5};
    assign wire3968 = {4'd7, 4'd6};
    assign wire3969 = {4'd7, 4'd6};
    assign wire3970 = {4'd7, 4'd6};
    assign wire3971 = {4'd7, 4'd6};
    assign wire3972 = {4'd7, 4'd6};
    assign wire3973 = {4'd9, 4'd8};
    assign wire3974 = {4'd7, 4'd6};
    assign wire3975 = {4'd7, 4'd6};
    assign wire3976 = {4'd8, 4'd7};
    assign wire3977 = {4'd8, 4'd7};
    assign wire3978 = {4'd8, 4'd7};
    assign wire3979 = {4'd8, 4'd7};
    assign wire3980 = {4'd8, 4'd7};
    assign wire3981 = {4'd8, 4'd7};
    assign wire3982 = {4'd8, 4'd7};
    assign wire3983 = {4'd8, 4'd7};
    assign wire3984 = {4'd9, 4'd8};
    assign wire3985 = {4'd9, 4'd8};
    assign wire3986 = {4'd9, 4'd8};
    assign wire3987 = {4'd9, 4'd8};
    assign wire3988 = {4'd9, 4'd8};
    assign wire3989 = {4'd9, 4'd8};
    assign wire3990 = {4'd9, 4'd8};
    assign wire3991 = {4'd9, 4'd8};
    assign wire3992 = {4'd7, 4'd6};
    assign wire3993 = {4'd7, 4'd6};
    assign wire3994 = {4'd7, 4'd6};
    assign wire3995 = {4'd7, 4'd6};
    assign wire3996 = {4'd7, 4'd6};
    assign wire3997 = {4'd7, 4'd6};
    assign wire3998 = {4'd7, 4'd6};
    assign wire3999 = {4'd7, 4'd6};
    assign wire4000 = {4'd8, 4'd6};
    assign wire4001 = {4'd8, 4'd6};
    assign wire4002 = {4'd8, 4'd6};
    assign wire4003 = {4'd8, 4'd6};
    assign wire4004 = {4'd8, 4'd6};
    assign wire4005 = {4'd10, 4'd8};
    assign wire4006 = {4'd8, 4'd6};
    assign wire4007 = {4'd8, 4'd6};
    assign wire4008 = {4'd9, 4'd7};
    assign wire4009 = {4'd9, 4'd7};
    assign wire4010 = {4'd9, 4'd7};
    assign wire4011 = {4'd9, 4'd7};
    assign wire4012 = {4'd9, 4'd7};
    assign wire4013 = {4'd9, 4'd7};
    assign wire4014 = {4'd9, 4'd7};
    assign wire4015 = {4'd9, 4'd7};
    assign wire4016 = {4'd10, 4'd8};
    assign wire4017 = {4'd10, 4'd8};
    assign wire4018 = {4'd10, 4'd8};
    assign wire4019 = {4'd10, 4'd8};
    assign wire4020 = {4'd10, 4'd8};
    assign wire4021 = {4'd10, 4'd8};
    assign wire4022 = {4'd10, 4'd8};
    assign wire4023 = {4'd10, 4'd8};
    assign wire4024 = {4'd8, 4'd6};
    assign wire4025 = {4'd8, 4'd6};
    assign wire4026 = {4'd8, 4'd6};
    assign wire4027 = {4'd8, 4'd6};
    assign wire4028 = {4'd8, 4'd6};
    assign wire4029 = {4'd8, 4'd6};
    assign wire4030 = {4'd8, 4'd6};
    assign wire4031 = {4'd8, 4'd6};
    assign wire4032 = {4'd10, 4'd6};
    assign wire4033 = {4'd10, 4'd6};
    assign wire4034 = {4'd10, 4'd6};
    assign wire4035 = {4'd10, 4'd6};
    assign wire4036 = {4'd10, 4'd6};
    assign wire4037 = {4'd12, 4'd8};
    assign wire4038 = {4'd10, 4'd6};
    assign wire4039 = {4'd10, 4'd6};
    assign wire4040 = {4'd11, 4'd7};
    assign wire4041 = {4'd11, 4'd7};
    assign wire4042 = {4'd11, 4'd7};
    assign wire4043 = {4'd11, 4'd7};
    assign wire4044 = {4'd11, 4'd7};
    assign wire4045 = {4'd11, 4'd7};
    assign wire4046 = {4'd11, 4'd7};
    assign wire4047 = {4'd11, 4'd7};
    assign wire4048 = {4'd12, 4'd8};
    assign wire4049 = {4'd12, 4'd8};
    assign wire4050 = {4'd12, 4'd8};
    assign wire4051 = {4'd12, 4'd8};
    assign wire4052 = {4'd12, 4'd8};
    assign wire4053 = {4'd12, 4'd8};
    assign wire4054 = {4'd12, 4'd8};
    assign wire4055 = {4'd12, 4'd8};
    assign wire4056 = {4'd10, 4'd6};
    assign wire4057 = {4'd10, 4'd6};
    assign wire4058 = {4'd10, 4'd6};
    assign wire4059 = {4'd10, 4'd6};
    assign wire4060 = {4'd10, 4'd6};
    assign wire4061 = {4'd10, 4'd6};
    assign wire4062 = {4'd10, 4'd6};
    assign wire4063 = {4'd10, 4'd6};
    assign wire4064 = {4'd12, 4'd6};
    assign wire4065 = {4'd12, 4'd6};
    assign wire4066 = {4'd12, 4'd6};
    assign wire4067 = {4'd12, 4'd6};
    assign wire4068 = {4'd12, 4'd6};
    assign wire4069 = {4'd14, 4'd8};
    assign wire4070 = {4'd12, 4'd6};
    assign wire4071 = {4'd12, 4'd6};
    assign wire4072 = {4'd13, 4'd7};
    assign wire4073 = {4'd13, 4'd7};
    assign wire4074 = {4'd13, 4'd7};
    assign wire4075 = {4'd13, 4'd7};
    assign wire4076 = {4'd13, 4'd7};
    assign wire4077 = {4'd13, 4'd7};
    assign wire4078 = {4'd13, 4'd7};
    assign wire4079 = {4'd13, 4'd7};
    assign wire4080 = {4'd14, 4'd8};
    assign wire4081 = {4'd14, 4'd8};
    assign wire4082 = {4'd14, 4'd8};
    assign wire4083 = {4'd14, 4'd8};
    assign wire4084 = {4'd14, 4'd8};
    assign wire4085 = {4'd14, 4'd8};
    assign wire4086 = {4'd14, 4'd8};
    assign wire4087 = {4'd14, 4'd8};
    assign wire4088 = {4'd12, 4'd6};
    assign wire4089 = {4'd12, 4'd6};
    assign wire4090 = {4'd12, 4'd6};
    assign wire4091 = {4'd12, 4'd6};
    assign wire4092 = {4'd12, 4'd6};
    assign wire4093 = {4'd12, 4'd6};
    assign wire4094 = {4'd12, 4'd6};
    assign wire4095 = {4'd12, 4'd6};


    equaln #(12) e0(.a(buffered_input), .b(12'b000000000000), .eq(weq0));
    equaln #(12) e1(.a(buffered_input), .b(12'b000000000001), .eq(weq1));
    equaln #(12) e2(.a(buffered_input), .b(12'b000000000010), .eq(weq2));
    equaln #(12) e3(.a(buffered_input), .b(12'b000000000011), .eq(weq3));
    equaln #(12) e4(.a(buffered_input), .b(12'b000000000100), .eq(weq4));
    equaln #(12) e5(.a(buffered_input), .b(12'b000000000101), .eq(weq5));
    equaln #(12) e6(.a(buffered_input), .b(12'b000000000110), .eq(weq6));
    equaln #(12) e7(.a(buffered_input), .b(12'b000000000111), .eq(weq7));
    equaln #(12) e8(.a(buffered_input), .b(12'b000000001000), .eq(weq8));
    equaln #(12) e9(.a(buffered_input), .b(12'b000000001001), .eq(weq9));
    equaln #(12) e10(.a(buffered_input), .b(12'b000000001010), .eq(weq10));
    equaln #(12) e11(.a(buffered_input), .b(12'b000000001011), .eq(weq11));
    equaln #(12) e12(.a(buffered_input), .b(12'b000000001100), .eq(weq12));
    equaln #(12) e13(.a(buffered_input), .b(12'b000000001101), .eq(weq13));
    equaln #(12) e14(.a(buffered_input), .b(12'b000000001110), .eq(weq14));
    equaln #(12) e15(.a(buffered_input), .b(12'b000000001111), .eq(weq15));
    equaln #(12) e16(.a(buffered_input), .b(12'b000000010000), .eq(weq16));
    equaln #(12) e17(.a(buffered_input), .b(12'b000000010001), .eq(weq17));
    equaln #(12) e18(.a(buffered_input), .b(12'b000000010010), .eq(weq18));
    equaln #(12) e19(.a(buffered_input), .b(12'b000000010011), .eq(weq19));
    equaln #(12) e20(.a(buffered_input), .b(12'b000000010100), .eq(weq20));
    equaln #(12) e21(.a(buffered_input), .b(12'b000000010101), .eq(weq21));
    equaln #(12) e22(.a(buffered_input), .b(12'b000000010110), .eq(weq22));
    equaln #(12) e23(.a(buffered_input), .b(12'b000000010111), .eq(weq23));
    equaln #(12) e24(.a(buffered_input), .b(12'b000000011000), .eq(weq24));
    equaln #(12) e25(.a(buffered_input), .b(12'b000000011001), .eq(weq25));
    equaln #(12) e26(.a(buffered_input), .b(12'b000000011010), .eq(weq26));
    equaln #(12) e27(.a(buffered_input), .b(12'b000000011011), .eq(weq27));
    equaln #(12) e28(.a(buffered_input), .b(12'b000000011100), .eq(weq28));
    equaln #(12) e29(.a(buffered_input), .b(12'b000000011101), .eq(weq29));
    equaln #(12) e30(.a(buffered_input), .b(12'b000000011110), .eq(weq30));
    equaln #(12) e31(.a(buffered_input), .b(12'b000000011111), .eq(weq31));
    equaln #(12) e32(.a(buffered_input), .b(12'b000000100000), .eq(weq32));
    equaln #(12) e33(.a(buffered_input), .b(12'b000000100001), .eq(weq33));
    equaln #(12) e34(.a(buffered_input), .b(12'b000000100010), .eq(weq34));
    equaln #(12) e35(.a(buffered_input), .b(12'b000000100011), .eq(weq35));
    equaln #(12) e36(.a(buffered_input), .b(12'b000000100100), .eq(weq36));
    equaln #(12) e37(.a(buffered_input), .b(12'b000000100101), .eq(weq37));
    equaln #(12) e38(.a(buffered_input), .b(12'b000000100110), .eq(weq38));
    equaln #(12) e39(.a(buffered_input), .b(12'b000000100111), .eq(weq39));
    equaln #(12) e40(.a(buffered_input), .b(12'b000000101000), .eq(weq40));
    equaln #(12) e41(.a(buffered_input), .b(12'b000000101001), .eq(weq41));
    equaln #(12) e42(.a(buffered_input), .b(12'b000000101010), .eq(weq42));
    equaln #(12) e43(.a(buffered_input), .b(12'b000000101011), .eq(weq43));
    equaln #(12) e44(.a(buffered_input), .b(12'b000000101100), .eq(weq44));
    equaln #(12) e45(.a(buffered_input), .b(12'b000000101101), .eq(weq45));
    equaln #(12) e46(.a(buffered_input), .b(12'b000000101110), .eq(weq46));
    equaln #(12) e47(.a(buffered_input), .b(12'b000000101111), .eq(weq47));
    equaln #(12) e48(.a(buffered_input), .b(12'b000000110000), .eq(weq48));
    equaln #(12) e49(.a(buffered_input), .b(12'b000000110001), .eq(weq49));
    equaln #(12) e50(.a(buffered_input), .b(12'b000000110010), .eq(weq50));
    equaln #(12) e51(.a(buffered_input), .b(12'b000000110011), .eq(weq51));
    equaln #(12) e52(.a(buffered_input), .b(12'b000000110100), .eq(weq52));
    equaln #(12) e53(.a(buffered_input), .b(12'b000000110101), .eq(weq53));
    equaln #(12) e54(.a(buffered_input), .b(12'b000000110110), .eq(weq54));
    equaln #(12) e55(.a(buffered_input), .b(12'b000000110111), .eq(weq55));
    equaln #(12) e56(.a(buffered_input), .b(12'b000000111000), .eq(weq56));
    equaln #(12) e57(.a(buffered_input), .b(12'b000000111001), .eq(weq57));
    equaln #(12) e58(.a(buffered_input), .b(12'b000000111010), .eq(weq58));
    equaln #(12) e59(.a(buffered_input), .b(12'b000000111011), .eq(weq59));
    equaln #(12) e60(.a(buffered_input), .b(12'b000000111100), .eq(weq60));
    equaln #(12) e61(.a(buffered_input), .b(12'b000000111101), .eq(weq61));
    equaln #(12) e62(.a(buffered_input), .b(12'b000000111110), .eq(weq62));
    equaln #(12) e63(.a(buffered_input), .b(12'b000000111111), .eq(weq63));
    equaln #(12) e64(.a(buffered_input), .b(12'b000001000000), .eq(weq64));
    equaln #(12) e65(.a(buffered_input), .b(12'b000001000001), .eq(weq65));
    equaln #(12) e66(.a(buffered_input), .b(12'b000001000010), .eq(weq66));
    equaln #(12) e67(.a(buffered_input), .b(12'b000001000011), .eq(weq67));
    equaln #(12) e68(.a(buffered_input), .b(12'b000001000100), .eq(weq68));
    equaln #(12) e69(.a(buffered_input), .b(12'b000001000101), .eq(weq69));
    equaln #(12) e70(.a(buffered_input), .b(12'b000001000110), .eq(weq70));
    equaln #(12) e71(.a(buffered_input), .b(12'b000001000111), .eq(weq71));
    equaln #(12) e72(.a(buffered_input), .b(12'b000001001000), .eq(weq72));
    equaln #(12) e73(.a(buffered_input), .b(12'b000001001001), .eq(weq73));
    equaln #(12) e74(.a(buffered_input), .b(12'b000001001010), .eq(weq74));
    equaln #(12) e75(.a(buffered_input), .b(12'b000001001011), .eq(weq75));
    equaln #(12) e76(.a(buffered_input), .b(12'b000001001100), .eq(weq76));
    equaln #(12) e77(.a(buffered_input), .b(12'b000001001101), .eq(weq77));
    equaln #(12) e78(.a(buffered_input), .b(12'b000001001110), .eq(weq78));
    equaln #(12) e79(.a(buffered_input), .b(12'b000001001111), .eq(weq79));
    equaln #(12) e80(.a(buffered_input), .b(12'b000001010000), .eq(weq80));
    equaln #(12) e81(.a(buffered_input), .b(12'b000001010001), .eq(weq81));
    equaln #(12) e82(.a(buffered_input), .b(12'b000001010010), .eq(weq82));
    equaln #(12) e83(.a(buffered_input), .b(12'b000001010011), .eq(weq83));
    equaln #(12) e84(.a(buffered_input), .b(12'b000001010100), .eq(weq84));
    equaln #(12) e85(.a(buffered_input), .b(12'b000001010101), .eq(weq85));
    equaln #(12) e86(.a(buffered_input), .b(12'b000001010110), .eq(weq86));
    equaln #(12) e87(.a(buffered_input), .b(12'b000001010111), .eq(weq87));
    equaln #(12) e88(.a(buffered_input), .b(12'b000001011000), .eq(weq88));
    equaln #(12) e89(.a(buffered_input), .b(12'b000001011001), .eq(weq89));
    equaln #(12) e90(.a(buffered_input), .b(12'b000001011010), .eq(weq90));
    equaln #(12) e91(.a(buffered_input), .b(12'b000001011011), .eq(weq91));
    equaln #(12) e92(.a(buffered_input), .b(12'b000001011100), .eq(weq92));
    equaln #(12) e93(.a(buffered_input), .b(12'b000001011101), .eq(weq93));
    equaln #(12) e94(.a(buffered_input), .b(12'b000001011110), .eq(weq94));
    equaln #(12) e95(.a(buffered_input), .b(12'b000001011111), .eq(weq95));
    equaln #(12) e96(.a(buffered_input), .b(12'b000001100000), .eq(weq96));
    equaln #(12) e97(.a(buffered_input), .b(12'b000001100001), .eq(weq97));
    equaln #(12) e98(.a(buffered_input), .b(12'b000001100010), .eq(weq98));
    equaln #(12) e99(.a(buffered_input), .b(12'b000001100011), .eq(weq99));
    equaln #(12) e100(.a(buffered_input), .b(12'b000001100100), .eq(weq100));
    equaln #(12) e101(.a(buffered_input), .b(12'b000001100101), .eq(weq101));
    equaln #(12) e102(.a(buffered_input), .b(12'b000001100110), .eq(weq102));
    equaln #(12) e103(.a(buffered_input), .b(12'b000001100111), .eq(weq103));
    equaln #(12) e104(.a(buffered_input), .b(12'b000001101000), .eq(weq104));
    equaln #(12) e105(.a(buffered_input), .b(12'b000001101001), .eq(weq105));
    equaln #(12) e106(.a(buffered_input), .b(12'b000001101010), .eq(weq106));
    equaln #(12) e107(.a(buffered_input), .b(12'b000001101011), .eq(weq107));
    equaln #(12) e108(.a(buffered_input), .b(12'b000001101100), .eq(weq108));
    equaln #(12) e109(.a(buffered_input), .b(12'b000001101101), .eq(weq109));
    equaln #(12) e110(.a(buffered_input), .b(12'b000001101110), .eq(weq110));
    equaln #(12) e111(.a(buffered_input), .b(12'b000001101111), .eq(weq111));
    equaln #(12) e112(.a(buffered_input), .b(12'b000001110000), .eq(weq112));
    equaln #(12) e113(.a(buffered_input), .b(12'b000001110001), .eq(weq113));
    equaln #(12) e114(.a(buffered_input), .b(12'b000001110010), .eq(weq114));
    equaln #(12) e115(.a(buffered_input), .b(12'b000001110011), .eq(weq115));
    equaln #(12) e116(.a(buffered_input), .b(12'b000001110100), .eq(weq116));
    equaln #(12) e117(.a(buffered_input), .b(12'b000001110101), .eq(weq117));
    equaln #(12) e118(.a(buffered_input), .b(12'b000001110110), .eq(weq118));
    equaln #(12) e119(.a(buffered_input), .b(12'b000001110111), .eq(weq119));
    equaln #(12) e120(.a(buffered_input), .b(12'b000001111000), .eq(weq120));
    equaln #(12) e121(.a(buffered_input), .b(12'b000001111001), .eq(weq121));
    equaln #(12) e122(.a(buffered_input), .b(12'b000001111010), .eq(weq122));
    equaln #(12) e123(.a(buffered_input), .b(12'b000001111011), .eq(weq123));
    equaln #(12) e124(.a(buffered_input), .b(12'b000001111100), .eq(weq124));
    equaln #(12) e125(.a(buffered_input), .b(12'b000001111101), .eq(weq125));
    equaln #(12) e126(.a(buffered_input), .b(12'b000001111110), .eq(weq126));
    equaln #(12) e127(.a(buffered_input), .b(12'b000001111111), .eq(weq127));
    equaln #(12) e128(.a(buffered_input), .b(12'b000010000000), .eq(weq128));
    equaln #(12) e129(.a(buffered_input), .b(12'b000010000001), .eq(weq129));
    equaln #(12) e130(.a(buffered_input), .b(12'b000010000010), .eq(weq130));
    equaln #(12) e131(.a(buffered_input), .b(12'b000010000011), .eq(weq131));
    equaln #(12) e132(.a(buffered_input), .b(12'b000010000100), .eq(weq132));
    equaln #(12) e133(.a(buffered_input), .b(12'b000010000101), .eq(weq133));
    equaln #(12) e134(.a(buffered_input), .b(12'b000010000110), .eq(weq134));
    equaln #(12) e135(.a(buffered_input), .b(12'b000010000111), .eq(weq135));
    equaln #(12) e136(.a(buffered_input), .b(12'b000010001000), .eq(weq136));
    equaln #(12) e137(.a(buffered_input), .b(12'b000010001001), .eq(weq137));
    equaln #(12) e138(.a(buffered_input), .b(12'b000010001010), .eq(weq138));
    equaln #(12) e139(.a(buffered_input), .b(12'b000010001011), .eq(weq139));
    equaln #(12) e140(.a(buffered_input), .b(12'b000010001100), .eq(weq140));
    equaln #(12) e141(.a(buffered_input), .b(12'b000010001101), .eq(weq141));
    equaln #(12) e142(.a(buffered_input), .b(12'b000010001110), .eq(weq142));
    equaln #(12) e143(.a(buffered_input), .b(12'b000010001111), .eq(weq143));
    equaln #(12) e144(.a(buffered_input), .b(12'b000010010000), .eq(weq144));
    equaln #(12) e145(.a(buffered_input), .b(12'b000010010001), .eq(weq145));
    equaln #(12) e146(.a(buffered_input), .b(12'b000010010010), .eq(weq146));
    equaln #(12) e147(.a(buffered_input), .b(12'b000010010011), .eq(weq147));
    equaln #(12) e148(.a(buffered_input), .b(12'b000010010100), .eq(weq148));
    equaln #(12) e149(.a(buffered_input), .b(12'b000010010101), .eq(weq149));
    equaln #(12) e150(.a(buffered_input), .b(12'b000010010110), .eq(weq150));
    equaln #(12) e151(.a(buffered_input), .b(12'b000010010111), .eq(weq151));
    equaln #(12) e152(.a(buffered_input), .b(12'b000010011000), .eq(weq152));
    equaln #(12) e153(.a(buffered_input), .b(12'b000010011001), .eq(weq153));
    equaln #(12) e154(.a(buffered_input), .b(12'b000010011010), .eq(weq154));
    equaln #(12) e155(.a(buffered_input), .b(12'b000010011011), .eq(weq155));
    equaln #(12) e156(.a(buffered_input), .b(12'b000010011100), .eq(weq156));
    equaln #(12) e157(.a(buffered_input), .b(12'b000010011101), .eq(weq157));
    equaln #(12) e158(.a(buffered_input), .b(12'b000010011110), .eq(weq158));
    equaln #(12) e159(.a(buffered_input), .b(12'b000010011111), .eq(weq159));
    equaln #(12) e160(.a(buffered_input), .b(12'b000010100000), .eq(weq160));
    equaln #(12) e161(.a(buffered_input), .b(12'b000010100001), .eq(weq161));
    equaln #(12) e162(.a(buffered_input), .b(12'b000010100010), .eq(weq162));
    equaln #(12) e163(.a(buffered_input), .b(12'b000010100011), .eq(weq163));
    equaln #(12) e164(.a(buffered_input), .b(12'b000010100100), .eq(weq164));
    equaln #(12) e165(.a(buffered_input), .b(12'b000010100101), .eq(weq165));
    equaln #(12) e166(.a(buffered_input), .b(12'b000010100110), .eq(weq166));
    equaln #(12) e167(.a(buffered_input), .b(12'b000010100111), .eq(weq167));
    equaln #(12) e168(.a(buffered_input), .b(12'b000010101000), .eq(weq168));
    equaln #(12) e169(.a(buffered_input), .b(12'b000010101001), .eq(weq169));
    equaln #(12) e170(.a(buffered_input), .b(12'b000010101010), .eq(weq170));
    equaln #(12) e171(.a(buffered_input), .b(12'b000010101011), .eq(weq171));
    equaln #(12) e172(.a(buffered_input), .b(12'b000010101100), .eq(weq172));
    equaln #(12) e173(.a(buffered_input), .b(12'b000010101101), .eq(weq173));
    equaln #(12) e174(.a(buffered_input), .b(12'b000010101110), .eq(weq174));
    equaln #(12) e175(.a(buffered_input), .b(12'b000010101111), .eq(weq175));
    equaln #(12) e176(.a(buffered_input), .b(12'b000010110000), .eq(weq176));
    equaln #(12) e177(.a(buffered_input), .b(12'b000010110001), .eq(weq177));
    equaln #(12) e178(.a(buffered_input), .b(12'b000010110010), .eq(weq178));
    equaln #(12) e179(.a(buffered_input), .b(12'b000010110011), .eq(weq179));
    equaln #(12) e180(.a(buffered_input), .b(12'b000010110100), .eq(weq180));
    equaln #(12) e181(.a(buffered_input), .b(12'b000010110101), .eq(weq181));
    equaln #(12) e182(.a(buffered_input), .b(12'b000010110110), .eq(weq182));
    equaln #(12) e183(.a(buffered_input), .b(12'b000010110111), .eq(weq183));
    equaln #(12) e184(.a(buffered_input), .b(12'b000010111000), .eq(weq184));
    equaln #(12) e185(.a(buffered_input), .b(12'b000010111001), .eq(weq185));
    equaln #(12) e186(.a(buffered_input), .b(12'b000010111010), .eq(weq186));
    equaln #(12) e187(.a(buffered_input), .b(12'b000010111011), .eq(weq187));
    equaln #(12) e188(.a(buffered_input), .b(12'b000010111100), .eq(weq188));
    equaln #(12) e189(.a(buffered_input), .b(12'b000010111101), .eq(weq189));
    equaln #(12) e190(.a(buffered_input), .b(12'b000010111110), .eq(weq190));
    equaln #(12) e191(.a(buffered_input), .b(12'b000010111111), .eq(weq191));
    equaln #(12) e192(.a(buffered_input), .b(12'b000011000000), .eq(weq192));
    equaln #(12) e193(.a(buffered_input), .b(12'b000011000001), .eq(weq193));
    equaln #(12) e194(.a(buffered_input), .b(12'b000011000010), .eq(weq194));
    equaln #(12) e195(.a(buffered_input), .b(12'b000011000011), .eq(weq195));
    equaln #(12) e196(.a(buffered_input), .b(12'b000011000100), .eq(weq196));
    equaln #(12) e197(.a(buffered_input), .b(12'b000011000101), .eq(weq197));
    equaln #(12) e198(.a(buffered_input), .b(12'b000011000110), .eq(weq198));
    equaln #(12) e199(.a(buffered_input), .b(12'b000011000111), .eq(weq199));
    equaln #(12) e200(.a(buffered_input), .b(12'b000011001000), .eq(weq200));
    equaln #(12) e201(.a(buffered_input), .b(12'b000011001001), .eq(weq201));
    equaln #(12) e202(.a(buffered_input), .b(12'b000011001010), .eq(weq202));
    equaln #(12) e203(.a(buffered_input), .b(12'b000011001011), .eq(weq203));
    equaln #(12) e204(.a(buffered_input), .b(12'b000011001100), .eq(weq204));
    equaln #(12) e205(.a(buffered_input), .b(12'b000011001101), .eq(weq205));
    equaln #(12) e206(.a(buffered_input), .b(12'b000011001110), .eq(weq206));
    equaln #(12) e207(.a(buffered_input), .b(12'b000011001111), .eq(weq207));
    equaln #(12) e208(.a(buffered_input), .b(12'b000011010000), .eq(weq208));
    equaln #(12) e209(.a(buffered_input), .b(12'b000011010001), .eq(weq209));
    equaln #(12) e210(.a(buffered_input), .b(12'b000011010010), .eq(weq210));
    equaln #(12) e211(.a(buffered_input), .b(12'b000011010011), .eq(weq211));
    equaln #(12) e212(.a(buffered_input), .b(12'b000011010100), .eq(weq212));
    equaln #(12) e213(.a(buffered_input), .b(12'b000011010101), .eq(weq213));
    equaln #(12) e214(.a(buffered_input), .b(12'b000011010110), .eq(weq214));
    equaln #(12) e215(.a(buffered_input), .b(12'b000011010111), .eq(weq215));
    equaln #(12) e216(.a(buffered_input), .b(12'b000011011000), .eq(weq216));
    equaln #(12) e217(.a(buffered_input), .b(12'b000011011001), .eq(weq217));
    equaln #(12) e218(.a(buffered_input), .b(12'b000011011010), .eq(weq218));
    equaln #(12) e219(.a(buffered_input), .b(12'b000011011011), .eq(weq219));
    equaln #(12) e220(.a(buffered_input), .b(12'b000011011100), .eq(weq220));
    equaln #(12) e221(.a(buffered_input), .b(12'b000011011101), .eq(weq221));
    equaln #(12) e222(.a(buffered_input), .b(12'b000011011110), .eq(weq222));
    equaln #(12) e223(.a(buffered_input), .b(12'b000011011111), .eq(weq223));
    equaln #(12) e224(.a(buffered_input), .b(12'b000011100000), .eq(weq224));
    equaln #(12) e225(.a(buffered_input), .b(12'b000011100001), .eq(weq225));
    equaln #(12) e226(.a(buffered_input), .b(12'b000011100010), .eq(weq226));
    equaln #(12) e227(.a(buffered_input), .b(12'b000011100011), .eq(weq227));
    equaln #(12) e228(.a(buffered_input), .b(12'b000011100100), .eq(weq228));
    equaln #(12) e229(.a(buffered_input), .b(12'b000011100101), .eq(weq229));
    equaln #(12) e230(.a(buffered_input), .b(12'b000011100110), .eq(weq230));
    equaln #(12) e231(.a(buffered_input), .b(12'b000011100111), .eq(weq231));
    equaln #(12) e232(.a(buffered_input), .b(12'b000011101000), .eq(weq232));
    equaln #(12) e233(.a(buffered_input), .b(12'b000011101001), .eq(weq233));
    equaln #(12) e234(.a(buffered_input), .b(12'b000011101010), .eq(weq234));
    equaln #(12) e235(.a(buffered_input), .b(12'b000011101011), .eq(weq235));
    equaln #(12) e236(.a(buffered_input), .b(12'b000011101100), .eq(weq236));
    equaln #(12) e237(.a(buffered_input), .b(12'b000011101101), .eq(weq237));
    equaln #(12) e238(.a(buffered_input), .b(12'b000011101110), .eq(weq238));
    equaln #(12) e239(.a(buffered_input), .b(12'b000011101111), .eq(weq239));
    equaln #(12) e240(.a(buffered_input), .b(12'b000011110000), .eq(weq240));
    equaln #(12) e241(.a(buffered_input), .b(12'b000011110001), .eq(weq241));
    equaln #(12) e242(.a(buffered_input), .b(12'b000011110010), .eq(weq242));
    equaln #(12) e243(.a(buffered_input), .b(12'b000011110011), .eq(weq243));
    equaln #(12) e244(.a(buffered_input), .b(12'b000011110100), .eq(weq244));
    equaln #(12) e245(.a(buffered_input), .b(12'b000011110101), .eq(weq245));
    equaln #(12) e246(.a(buffered_input), .b(12'b000011110110), .eq(weq246));
    equaln #(12) e247(.a(buffered_input), .b(12'b000011110111), .eq(weq247));
    equaln #(12) e248(.a(buffered_input), .b(12'b000011111000), .eq(weq248));
    equaln #(12) e249(.a(buffered_input), .b(12'b000011111001), .eq(weq249));
    equaln #(12) e250(.a(buffered_input), .b(12'b000011111010), .eq(weq250));
    equaln #(12) e251(.a(buffered_input), .b(12'b000011111011), .eq(weq251));
    equaln #(12) e252(.a(buffered_input), .b(12'b000011111100), .eq(weq252));
    equaln #(12) e253(.a(buffered_input), .b(12'b000011111101), .eq(weq253));
    equaln #(12) e254(.a(buffered_input), .b(12'b000011111110), .eq(weq254));
    equaln #(12) e255(.a(buffered_input), .b(12'b000011111111), .eq(weq255));
    equaln #(12) e256(.a(buffered_input), .b(12'b000100000000), .eq(weq256));
    equaln #(12) e257(.a(buffered_input), .b(12'b000100000001), .eq(weq257));
    equaln #(12) e258(.a(buffered_input), .b(12'b000100000010), .eq(weq258));
    equaln #(12) e259(.a(buffered_input), .b(12'b000100000011), .eq(weq259));
    equaln #(12) e260(.a(buffered_input), .b(12'b000100000100), .eq(weq260));
    equaln #(12) e261(.a(buffered_input), .b(12'b000100000101), .eq(weq261));
    equaln #(12) e262(.a(buffered_input), .b(12'b000100000110), .eq(weq262));
    equaln #(12) e263(.a(buffered_input), .b(12'b000100000111), .eq(weq263));
    equaln #(12) e264(.a(buffered_input), .b(12'b000100001000), .eq(weq264));
    equaln #(12) e265(.a(buffered_input), .b(12'b000100001001), .eq(weq265));
    equaln #(12) e266(.a(buffered_input), .b(12'b000100001010), .eq(weq266));
    equaln #(12) e267(.a(buffered_input), .b(12'b000100001011), .eq(weq267));
    equaln #(12) e268(.a(buffered_input), .b(12'b000100001100), .eq(weq268));
    equaln #(12) e269(.a(buffered_input), .b(12'b000100001101), .eq(weq269));
    equaln #(12) e270(.a(buffered_input), .b(12'b000100001110), .eq(weq270));
    equaln #(12) e271(.a(buffered_input), .b(12'b000100001111), .eq(weq271));
    equaln #(12) e272(.a(buffered_input), .b(12'b000100010000), .eq(weq272));
    equaln #(12) e273(.a(buffered_input), .b(12'b000100010001), .eq(weq273));
    equaln #(12) e274(.a(buffered_input), .b(12'b000100010010), .eq(weq274));
    equaln #(12) e275(.a(buffered_input), .b(12'b000100010011), .eq(weq275));
    equaln #(12) e276(.a(buffered_input), .b(12'b000100010100), .eq(weq276));
    equaln #(12) e277(.a(buffered_input), .b(12'b000100010101), .eq(weq277));
    equaln #(12) e278(.a(buffered_input), .b(12'b000100010110), .eq(weq278));
    equaln #(12) e279(.a(buffered_input), .b(12'b000100010111), .eq(weq279));
    equaln #(12) e280(.a(buffered_input), .b(12'b000100011000), .eq(weq280));
    equaln #(12) e281(.a(buffered_input), .b(12'b000100011001), .eq(weq281));
    equaln #(12) e282(.a(buffered_input), .b(12'b000100011010), .eq(weq282));
    equaln #(12) e283(.a(buffered_input), .b(12'b000100011011), .eq(weq283));
    equaln #(12) e284(.a(buffered_input), .b(12'b000100011100), .eq(weq284));
    equaln #(12) e285(.a(buffered_input), .b(12'b000100011101), .eq(weq285));
    equaln #(12) e286(.a(buffered_input), .b(12'b000100011110), .eq(weq286));
    equaln #(12) e287(.a(buffered_input), .b(12'b000100011111), .eq(weq287));
    equaln #(12) e288(.a(buffered_input), .b(12'b000100100000), .eq(weq288));
    equaln #(12) e289(.a(buffered_input), .b(12'b000100100001), .eq(weq289));
    equaln #(12) e290(.a(buffered_input), .b(12'b000100100010), .eq(weq290));
    equaln #(12) e291(.a(buffered_input), .b(12'b000100100011), .eq(weq291));
    equaln #(12) e292(.a(buffered_input), .b(12'b000100100100), .eq(weq292));
    equaln #(12) e293(.a(buffered_input), .b(12'b000100100101), .eq(weq293));
    equaln #(12) e294(.a(buffered_input), .b(12'b000100100110), .eq(weq294));
    equaln #(12) e295(.a(buffered_input), .b(12'b000100100111), .eq(weq295));
    equaln #(12) e296(.a(buffered_input), .b(12'b000100101000), .eq(weq296));
    equaln #(12) e297(.a(buffered_input), .b(12'b000100101001), .eq(weq297));
    equaln #(12) e298(.a(buffered_input), .b(12'b000100101010), .eq(weq298));
    equaln #(12) e299(.a(buffered_input), .b(12'b000100101011), .eq(weq299));
    equaln #(12) e300(.a(buffered_input), .b(12'b000100101100), .eq(weq300));
    equaln #(12) e301(.a(buffered_input), .b(12'b000100101101), .eq(weq301));
    equaln #(12) e302(.a(buffered_input), .b(12'b000100101110), .eq(weq302));
    equaln #(12) e303(.a(buffered_input), .b(12'b000100101111), .eq(weq303));
    equaln #(12) e304(.a(buffered_input), .b(12'b000100110000), .eq(weq304));
    equaln #(12) e305(.a(buffered_input), .b(12'b000100110001), .eq(weq305));
    equaln #(12) e306(.a(buffered_input), .b(12'b000100110010), .eq(weq306));
    equaln #(12) e307(.a(buffered_input), .b(12'b000100110011), .eq(weq307));
    equaln #(12) e308(.a(buffered_input), .b(12'b000100110100), .eq(weq308));
    equaln #(12) e309(.a(buffered_input), .b(12'b000100110101), .eq(weq309));
    equaln #(12) e310(.a(buffered_input), .b(12'b000100110110), .eq(weq310));
    equaln #(12) e311(.a(buffered_input), .b(12'b000100110111), .eq(weq311));
    equaln #(12) e312(.a(buffered_input), .b(12'b000100111000), .eq(weq312));
    equaln #(12) e313(.a(buffered_input), .b(12'b000100111001), .eq(weq313));
    equaln #(12) e314(.a(buffered_input), .b(12'b000100111010), .eq(weq314));
    equaln #(12) e315(.a(buffered_input), .b(12'b000100111011), .eq(weq315));
    equaln #(12) e316(.a(buffered_input), .b(12'b000100111100), .eq(weq316));
    equaln #(12) e317(.a(buffered_input), .b(12'b000100111101), .eq(weq317));
    equaln #(12) e318(.a(buffered_input), .b(12'b000100111110), .eq(weq318));
    equaln #(12) e319(.a(buffered_input), .b(12'b000100111111), .eq(weq319));
    equaln #(12) e320(.a(buffered_input), .b(12'b000101000000), .eq(weq320));
    equaln #(12) e321(.a(buffered_input), .b(12'b000101000001), .eq(weq321));
    equaln #(12) e322(.a(buffered_input), .b(12'b000101000010), .eq(weq322));
    equaln #(12) e323(.a(buffered_input), .b(12'b000101000011), .eq(weq323));
    equaln #(12) e324(.a(buffered_input), .b(12'b000101000100), .eq(weq324));
    equaln #(12) e325(.a(buffered_input), .b(12'b000101000101), .eq(weq325));
    equaln #(12) e326(.a(buffered_input), .b(12'b000101000110), .eq(weq326));
    equaln #(12) e327(.a(buffered_input), .b(12'b000101000111), .eq(weq327));
    equaln #(12) e328(.a(buffered_input), .b(12'b000101001000), .eq(weq328));
    equaln #(12) e329(.a(buffered_input), .b(12'b000101001001), .eq(weq329));
    equaln #(12) e330(.a(buffered_input), .b(12'b000101001010), .eq(weq330));
    equaln #(12) e331(.a(buffered_input), .b(12'b000101001011), .eq(weq331));
    equaln #(12) e332(.a(buffered_input), .b(12'b000101001100), .eq(weq332));
    equaln #(12) e333(.a(buffered_input), .b(12'b000101001101), .eq(weq333));
    equaln #(12) e334(.a(buffered_input), .b(12'b000101001110), .eq(weq334));
    equaln #(12) e335(.a(buffered_input), .b(12'b000101001111), .eq(weq335));
    equaln #(12) e336(.a(buffered_input), .b(12'b000101010000), .eq(weq336));
    equaln #(12) e337(.a(buffered_input), .b(12'b000101010001), .eq(weq337));
    equaln #(12) e338(.a(buffered_input), .b(12'b000101010010), .eq(weq338));
    equaln #(12) e339(.a(buffered_input), .b(12'b000101010011), .eq(weq339));
    equaln #(12) e340(.a(buffered_input), .b(12'b000101010100), .eq(weq340));
    equaln #(12) e341(.a(buffered_input), .b(12'b000101010101), .eq(weq341));
    equaln #(12) e342(.a(buffered_input), .b(12'b000101010110), .eq(weq342));
    equaln #(12) e343(.a(buffered_input), .b(12'b000101010111), .eq(weq343));
    equaln #(12) e344(.a(buffered_input), .b(12'b000101011000), .eq(weq344));
    equaln #(12) e345(.a(buffered_input), .b(12'b000101011001), .eq(weq345));
    equaln #(12) e346(.a(buffered_input), .b(12'b000101011010), .eq(weq346));
    equaln #(12) e347(.a(buffered_input), .b(12'b000101011011), .eq(weq347));
    equaln #(12) e348(.a(buffered_input), .b(12'b000101011100), .eq(weq348));
    equaln #(12) e349(.a(buffered_input), .b(12'b000101011101), .eq(weq349));
    equaln #(12) e350(.a(buffered_input), .b(12'b000101011110), .eq(weq350));
    equaln #(12) e351(.a(buffered_input), .b(12'b000101011111), .eq(weq351));
    equaln #(12) e352(.a(buffered_input), .b(12'b000101100000), .eq(weq352));
    equaln #(12) e353(.a(buffered_input), .b(12'b000101100001), .eq(weq353));
    equaln #(12) e354(.a(buffered_input), .b(12'b000101100010), .eq(weq354));
    equaln #(12) e355(.a(buffered_input), .b(12'b000101100011), .eq(weq355));
    equaln #(12) e356(.a(buffered_input), .b(12'b000101100100), .eq(weq356));
    equaln #(12) e357(.a(buffered_input), .b(12'b000101100101), .eq(weq357));
    equaln #(12) e358(.a(buffered_input), .b(12'b000101100110), .eq(weq358));
    equaln #(12) e359(.a(buffered_input), .b(12'b000101100111), .eq(weq359));
    equaln #(12) e360(.a(buffered_input), .b(12'b000101101000), .eq(weq360));
    equaln #(12) e361(.a(buffered_input), .b(12'b000101101001), .eq(weq361));
    equaln #(12) e362(.a(buffered_input), .b(12'b000101101010), .eq(weq362));
    equaln #(12) e363(.a(buffered_input), .b(12'b000101101011), .eq(weq363));
    equaln #(12) e364(.a(buffered_input), .b(12'b000101101100), .eq(weq364));
    equaln #(12) e365(.a(buffered_input), .b(12'b000101101101), .eq(weq365));
    equaln #(12) e366(.a(buffered_input), .b(12'b000101101110), .eq(weq366));
    equaln #(12) e367(.a(buffered_input), .b(12'b000101101111), .eq(weq367));
    equaln #(12) e368(.a(buffered_input), .b(12'b000101110000), .eq(weq368));
    equaln #(12) e369(.a(buffered_input), .b(12'b000101110001), .eq(weq369));
    equaln #(12) e370(.a(buffered_input), .b(12'b000101110010), .eq(weq370));
    equaln #(12) e371(.a(buffered_input), .b(12'b000101110011), .eq(weq371));
    equaln #(12) e372(.a(buffered_input), .b(12'b000101110100), .eq(weq372));
    equaln #(12) e373(.a(buffered_input), .b(12'b000101110101), .eq(weq373));
    equaln #(12) e374(.a(buffered_input), .b(12'b000101110110), .eq(weq374));
    equaln #(12) e375(.a(buffered_input), .b(12'b000101110111), .eq(weq375));
    equaln #(12) e376(.a(buffered_input), .b(12'b000101111000), .eq(weq376));
    equaln #(12) e377(.a(buffered_input), .b(12'b000101111001), .eq(weq377));
    equaln #(12) e378(.a(buffered_input), .b(12'b000101111010), .eq(weq378));
    equaln #(12) e379(.a(buffered_input), .b(12'b000101111011), .eq(weq379));
    equaln #(12) e380(.a(buffered_input), .b(12'b000101111100), .eq(weq380));
    equaln #(12) e381(.a(buffered_input), .b(12'b000101111101), .eq(weq381));
    equaln #(12) e382(.a(buffered_input), .b(12'b000101111110), .eq(weq382));
    equaln #(12) e383(.a(buffered_input), .b(12'b000101111111), .eq(weq383));
    equaln #(12) e384(.a(buffered_input), .b(12'b000110000000), .eq(weq384));
    equaln #(12) e385(.a(buffered_input), .b(12'b000110000001), .eq(weq385));
    equaln #(12) e386(.a(buffered_input), .b(12'b000110000010), .eq(weq386));
    equaln #(12) e387(.a(buffered_input), .b(12'b000110000011), .eq(weq387));
    equaln #(12) e388(.a(buffered_input), .b(12'b000110000100), .eq(weq388));
    equaln #(12) e389(.a(buffered_input), .b(12'b000110000101), .eq(weq389));
    equaln #(12) e390(.a(buffered_input), .b(12'b000110000110), .eq(weq390));
    equaln #(12) e391(.a(buffered_input), .b(12'b000110000111), .eq(weq391));
    equaln #(12) e392(.a(buffered_input), .b(12'b000110001000), .eq(weq392));
    equaln #(12) e393(.a(buffered_input), .b(12'b000110001001), .eq(weq393));
    equaln #(12) e394(.a(buffered_input), .b(12'b000110001010), .eq(weq394));
    equaln #(12) e395(.a(buffered_input), .b(12'b000110001011), .eq(weq395));
    equaln #(12) e396(.a(buffered_input), .b(12'b000110001100), .eq(weq396));
    equaln #(12) e397(.a(buffered_input), .b(12'b000110001101), .eq(weq397));
    equaln #(12) e398(.a(buffered_input), .b(12'b000110001110), .eq(weq398));
    equaln #(12) e399(.a(buffered_input), .b(12'b000110001111), .eq(weq399));
    equaln #(12) e400(.a(buffered_input), .b(12'b000110010000), .eq(weq400));
    equaln #(12) e401(.a(buffered_input), .b(12'b000110010001), .eq(weq401));
    equaln #(12) e402(.a(buffered_input), .b(12'b000110010010), .eq(weq402));
    equaln #(12) e403(.a(buffered_input), .b(12'b000110010011), .eq(weq403));
    equaln #(12) e404(.a(buffered_input), .b(12'b000110010100), .eq(weq404));
    equaln #(12) e405(.a(buffered_input), .b(12'b000110010101), .eq(weq405));
    equaln #(12) e406(.a(buffered_input), .b(12'b000110010110), .eq(weq406));
    equaln #(12) e407(.a(buffered_input), .b(12'b000110010111), .eq(weq407));
    equaln #(12) e408(.a(buffered_input), .b(12'b000110011000), .eq(weq408));
    equaln #(12) e409(.a(buffered_input), .b(12'b000110011001), .eq(weq409));
    equaln #(12) e410(.a(buffered_input), .b(12'b000110011010), .eq(weq410));
    equaln #(12) e411(.a(buffered_input), .b(12'b000110011011), .eq(weq411));
    equaln #(12) e412(.a(buffered_input), .b(12'b000110011100), .eq(weq412));
    equaln #(12) e413(.a(buffered_input), .b(12'b000110011101), .eq(weq413));
    equaln #(12) e414(.a(buffered_input), .b(12'b000110011110), .eq(weq414));
    equaln #(12) e415(.a(buffered_input), .b(12'b000110011111), .eq(weq415));
    equaln #(12) e416(.a(buffered_input), .b(12'b000110100000), .eq(weq416));
    equaln #(12) e417(.a(buffered_input), .b(12'b000110100001), .eq(weq417));
    equaln #(12) e418(.a(buffered_input), .b(12'b000110100010), .eq(weq418));
    equaln #(12) e419(.a(buffered_input), .b(12'b000110100011), .eq(weq419));
    equaln #(12) e420(.a(buffered_input), .b(12'b000110100100), .eq(weq420));
    equaln #(12) e421(.a(buffered_input), .b(12'b000110100101), .eq(weq421));
    equaln #(12) e422(.a(buffered_input), .b(12'b000110100110), .eq(weq422));
    equaln #(12) e423(.a(buffered_input), .b(12'b000110100111), .eq(weq423));
    equaln #(12) e424(.a(buffered_input), .b(12'b000110101000), .eq(weq424));
    equaln #(12) e425(.a(buffered_input), .b(12'b000110101001), .eq(weq425));
    equaln #(12) e426(.a(buffered_input), .b(12'b000110101010), .eq(weq426));
    equaln #(12) e427(.a(buffered_input), .b(12'b000110101011), .eq(weq427));
    equaln #(12) e428(.a(buffered_input), .b(12'b000110101100), .eq(weq428));
    equaln #(12) e429(.a(buffered_input), .b(12'b000110101101), .eq(weq429));
    equaln #(12) e430(.a(buffered_input), .b(12'b000110101110), .eq(weq430));
    equaln #(12) e431(.a(buffered_input), .b(12'b000110101111), .eq(weq431));
    equaln #(12) e432(.a(buffered_input), .b(12'b000110110000), .eq(weq432));
    equaln #(12) e433(.a(buffered_input), .b(12'b000110110001), .eq(weq433));
    equaln #(12) e434(.a(buffered_input), .b(12'b000110110010), .eq(weq434));
    equaln #(12) e435(.a(buffered_input), .b(12'b000110110011), .eq(weq435));
    equaln #(12) e436(.a(buffered_input), .b(12'b000110110100), .eq(weq436));
    equaln #(12) e437(.a(buffered_input), .b(12'b000110110101), .eq(weq437));
    equaln #(12) e438(.a(buffered_input), .b(12'b000110110110), .eq(weq438));
    equaln #(12) e439(.a(buffered_input), .b(12'b000110110111), .eq(weq439));
    equaln #(12) e440(.a(buffered_input), .b(12'b000110111000), .eq(weq440));
    equaln #(12) e441(.a(buffered_input), .b(12'b000110111001), .eq(weq441));
    equaln #(12) e442(.a(buffered_input), .b(12'b000110111010), .eq(weq442));
    equaln #(12) e443(.a(buffered_input), .b(12'b000110111011), .eq(weq443));
    equaln #(12) e444(.a(buffered_input), .b(12'b000110111100), .eq(weq444));
    equaln #(12) e445(.a(buffered_input), .b(12'b000110111101), .eq(weq445));
    equaln #(12) e446(.a(buffered_input), .b(12'b000110111110), .eq(weq446));
    equaln #(12) e447(.a(buffered_input), .b(12'b000110111111), .eq(weq447));
    equaln #(12) e448(.a(buffered_input), .b(12'b000111000000), .eq(weq448));
    equaln #(12) e449(.a(buffered_input), .b(12'b000111000001), .eq(weq449));
    equaln #(12) e450(.a(buffered_input), .b(12'b000111000010), .eq(weq450));
    equaln #(12) e451(.a(buffered_input), .b(12'b000111000011), .eq(weq451));
    equaln #(12) e452(.a(buffered_input), .b(12'b000111000100), .eq(weq452));
    equaln #(12) e453(.a(buffered_input), .b(12'b000111000101), .eq(weq453));
    equaln #(12) e454(.a(buffered_input), .b(12'b000111000110), .eq(weq454));
    equaln #(12) e455(.a(buffered_input), .b(12'b000111000111), .eq(weq455));
    equaln #(12) e456(.a(buffered_input), .b(12'b000111001000), .eq(weq456));
    equaln #(12) e457(.a(buffered_input), .b(12'b000111001001), .eq(weq457));
    equaln #(12) e458(.a(buffered_input), .b(12'b000111001010), .eq(weq458));
    equaln #(12) e459(.a(buffered_input), .b(12'b000111001011), .eq(weq459));
    equaln #(12) e460(.a(buffered_input), .b(12'b000111001100), .eq(weq460));
    equaln #(12) e461(.a(buffered_input), .b(12'b000111001101), .eq(weq461));
    equaln #(12) e462(.a(buffered_input), .b(12'b000111001110), .eq(weq462));
    equaln #(12) e463(.a(buffered_input), .b(12'b000111001111), .eq(weq463));
    equaln #(12) e464(.a(buffered_input), .b(12'b000111010000), .eq(weq464));
    equaln #(12) e465(.a(buffered_input), .b(12'b000111010001), .eq(weq465));
    equaln #(12) e466(.a(buffered_input), .b(12'b000111010010), .eq(weq466));
    equaln #(12) e467(.a(buffered_input), .b(12'b000111010011), .eq(weq467));
    equaln #(12) e468(.a(buffered_input), .b(12'b000111010100), .eq(weq468));
    equaln #(12) e469(.a(buffered_input), .b(12'b000111010101), .eq(weq469));
    equaln #(12) e470(.a(buffered_input), .b(12'b000111010110), .eq(weq470));
    equaln #(12) e471(.a(buffered_input), .b(12'b000111010111), .eq(weq471));
    equaln #(12) e472(.a(buffered_input), .b(12'b000111011000), .eq(weq472));
    equaln #(12) e473(.a(buffered_input), .b(12'b000111011001), .eq(weq473));
    equaln #(12) e474(.a(buffered_input), .b(12'b000111011010), .eq(weq474));
    equaln #(12) e475(.a(buffered_input), .b(12'b000111011011), .eq(weq475));
    equaln #(12) e476(.a(buffered_input), .b(12'b000111011100), .eq(weq476));
    equaln #(12) e477(.a(buffered_input), .b(12'b000111011101), .eq(weq477));
    equaln #(12) e478(.a(buffered_input), .b(12'b000111011110), .eq(weq478));
    equaln #(12) e479(.a(buffered_input), .b(12'b000111011111), .eq(weq479));
    equaln #(12) e480(.a(buffered_input), .b(12'b000111100000), .eq(weq480));
    equaln #(12) e481(.a(buffered_input), .b(12'b000111100001), .eq(weq481));
    equaln #(12) e482(.a(buffered_input), .b(12'b000111100010), .eq(weq482));
    equaln #(12) e483(.a(buffered_input), .b(12'b000111100011), .eq(weq483));
    equaln #(12) e484(.a(buffered_input), .b(12'b000111100100), .eq(weq484));
    equaln #(12) e485(.a(buffered_input), .b(12'b000111100101), .eq(weq485));
    equaln #(12) e486(.a(buffered_input), .b(12'b000111100110), .eq(weq486));
    equaln #(12) e487(.a(buffered_input), .b(12'b000111100111), .eq(weq487));
    equaln #(12) e488(.a(buffered_input), .b(12'b000111101000), .eq(weq488));
    equaln #(12) e489(.a(buffered_input), .b(12'b000111101001), .eq(weq489));
    equaln #(12) e490(.a(buffered_input), .b(12'b000111101010), .eq(weq490));
    equaln #(12) e491(.a(buffered_input), .b(12'b000111101011), .eq(weq491));
    equaln #(12) e492(.a(buffered_input), .b(12'b000111101100), .eq(weq492));
    equaln #(12) e493(.a(buffered_input), .b(12'b000111101101), .eq(weq493));
    equaln #(12) e494(.a(buffered_input), .b(12'b000111101110), .eq(weq494));
    equaln #(12) e495(.a(buffered_input), .b(12'b000111101111), .eq(weq495));
    equaln #(12) e496(.a(buffered_input), .b(12'b000111110000), .eq(weq496));
    equaln #(12) e497(.a(buffered_input), .b(12'b000111110001), .eq(weq497));
    equaln #(12) e498(.a(buffered_input), .b(12'b000111110010), .eq(weq498));
    equaln #(12) e499(.a(buffered_input), .b(12'b000111110011), .eq(weq499));
    equaln #(12) e500(.a(buffered_input), .b(12'b000111110100), .eq(weq500));
    equaln #(12) e501(.a(buffered_input), .b(12'b000111110101), .eq(weq501));
    equaln #(12) e502(.a(buffered_input), .b(12'b000111110110), .eq(weq502));
    equaln #(12) e503(.a(buffered_input), .b(12'b000111110111), .eq(weq503));
    equaln #(12) e504(.a(buffered_input), .b(12'b000111111000), .eq(weq504));
    equaln #(12) e505(.a(buffered_input), .b(12'b000111111001), .eq(weq505));
    equaln #(12) e506(.a(buffered_input), .b(12'b000111111010), .eq(weq506));
    equaln #(12) e507(.a(buffered_input), .b(12'b000111111011), .eq(weq507));
    equaln #(12) e508(.a(buffered_input), .b(12'b000111111100), .eq(weq508));
    equaln #(12) e509(.a(buffered_input), .b(12'b000111111101), .eq(weq509));
    equaln #(12) e510(.a(buffered_input), .b(12'b000111111110), .eq(weq510));
    equaln #(12) e511(.a(buffered_input), .b(12'b000111111111), .eq(weq511));
    equaln #(12) e512(.a(buffered_input), .b(12'b001000000000), .eq(weq512));
    equaln #(12) e513(.a(buffered_input), .b(12'b001000000001), .eq(weq513));
    equaln #(12) e514(.a(buffered_input), .b(12'b001000000010), .eq(weq514));
    equaln #(12) e515(.a(buffered_input), .b(12'b001000000011), .eq(weq515));
    equaln #(12) e516(.a(buffered_input), .b(12'b001000000100), .eq(weq516));
    equaln #(12) e517(.a(buffered_input), .b(12'b001000000101), .eq(weq517));
    equaln #(12) e518(.a(buffered_input), .b(12'b001000000110), .eq(weq518));
    equaln #(12) e519(.a(buffered_input), .b(12'b001000000111), .eq(weq519));
    equaln #(12) e520(.a(buffered_input), .b(12'b001000001000), .eq(weq520));
    equaln #(12) e521(.a(buffered_input), .b(12'b001000001001), .eq(weq521));
    equaln #(12) e522(.a(buffered_input), .b(12'b001000001010), .eq(weq522));
    equaln #(12) e523(.a(buffered_input), .b(12'b001000001011), .eq(weq523));
    equaln #(12) e524(.a(buffered_input), .b(12'b001000001100), .eq(weq524));
    equaln #(12) e525(.a(buffered_input), .b(12'b001000001101), .eq(weq525));
    equaln #(12) e526(.a(buffered_input), .b(12'b001000001110), .eq(weq526));
    equaln #(12) e527(.a(buffered_input), .b(12'b001000001111), .eq(weq527));
    equaln #(12) e528(.a(buffered_input), .b(12'b001000010000), .eq(weq528));
    equaln #(12) e529(.a(buffered_input), .b(12'b001000010001), .eq(weq529));
    equaln #(12) e530(.a(buffered_input), .b(12'b001000010010), .eq(weq530));
    equaln #(12) e531(.a(buffered_input), .b(12'b001000010011), .eq(weq531));
    equaln #(12) e532(.a(buffered_input), .b(12'b001000010100), .eq(weq532));
    equaln #(12) e533(.a(buffered_input), .b(12'b001000010101), .eq(weq533));
    equaln #(12) e534(.a(buffered_input), .b(12'b001000010110), .eq(weq534));
    equaln #(12) e535(.a(buffered_input), .b(12'b001000010111), .eq(weq535));
    equaln #(12) e536(.a(buffered_input), .b(12'b001000011000), .eq(weq536));
    equaln #(12) e537(.a(buffered_input), .b(12'b001000011001), .eq(weq537));
    equaln #(12) e538(.a(buffered_input), .b(12'b001000011010), .eq(weq538));
    equaln #(12) e539(.a(buffered_input), .b(12'b001000011011), .eq(weq539));
    equaln #(12) e540(.a(buffered_input), .b(12'b001000011100), .eq(weq540));
    equaln #(12) e541(.a(buffered_input), .b(12'b001000011101), .eq(weq541));
    equaln #(12) e542(.a(buffered_input), .b(12'b001000011110), .eq(weq542));
    equaln #(12) e543(.a(buffered_input), .b(12'b001000011111), .eq(weq543));
    equaln #(12) e544(.a(buffered_input), .b(12'b001000100000), .eq(weq544));
    equaln #(12) e545(.a(buffered_input), .b(12'b001000100001), .eq(weq545));
    equaln #(12) e546(.a(buffered_input), .b(12'b001000100010), .eq(weq546));
    equaln #(12) e547(.a(buffered_input), .b(12'b001000100011), .eq(weq547));
    equaln #(12) e548(.a(buffered_input), .b(12'b001000100100), .eq(weq548));
    equaln #(12) e549(.a(buffered_input), .b(12'b001000100101), .eq(weq549));
    equaln #(12) e550(.a(buffered_input), .b(12'b001000100110), .eq(weq550));
    equaln #(12) e551(.a(buffered_input), .b(12'b001000100111), .eq(weq551));
    equaln #(12) e552(.a(buffered_input), .b(12'b001000101000), .eq(weq552));
    equaln #(12) e553(.a(buffered_input), .b(12'b001000101001), .eq(weq553));
    equaln #(12) e554(.a(buffered_input), .b(12'b001000101010), .eq(weq554));
    equaln #(12) e555(.a(buffered_input), .b(12'b001000101011), .eq(weq555));
    equaln #(12) e556(.a(buffered_input), .b(12'b001000101100), .eq(weq556));
    equaln #(12) e557(.a(buffered_input), .b(12'b001000101101), .eq(weq557));
    equaln #(12) e558(.a(buffered_input), .b(12'b001000101110), .eq(weq558));
    equaln #(12) e559(.a(buffered_input), .b(12'b001000101111), .eq(weq559));
    equaln #(12) e560(.a(buffered_input), .b(12'b001000110000), .eq(weq560));
    equaln #(12) e561(.a(buffered_input), .b(12'b001000110001), .eq(weq561));
    equaln #(12) e562(.a(buffered_input), .b(12'b001000110010), .eq(weq562));
    equaln #(12) e563(.a(buffered_input), .b(12'b001000110011), .eq(weq563));
    equaln #(12) e564(.a(buffered_input), .b(12'b001000110100), .eq(weq564));
    equaln #(12) e565(.a(buffered_input), .b(12'b001000110101), .eq(weq565));
    equaln #(12) e566(.a(buffered_input), .b(12'b001000110110), .eq(weq566));
    equaln #(12) e567(.a(buffered_input), .b(12'b001000110111), .eq(weq567));
    equaln #(12) e568(.a(buffered_input), .b(12'b001000111000), .eq(weq568));
    equaln #(12) e569(.a(buffered_input), .b(12'b001000111001), .eq(weq569));
    equaln #(12) e570(.a(buffered_input), .b(12'b001000111010), .eq(weq570));
    equaln #(12) e571(.a(buffered_input), .b(12'b001000111011), .eq(weq571));
    equaln #(12) e572(.a(buffered_input), .b(12'b001000111100), .eq(weq572));
    equaln #(12) e573(.a(buffered_input), .b(12'b001000111101), .eq(weq573));
    equaln #(12) e574(.a(buffered_input), .b(12'b001000111110), .eq(weq574));
    equaln #(12) e575(.a(buffered_input), .b(12'b001000111111), .eq(weq575));
    equaln #(12) e576(.a(buffered_input), .b(12'b001001000000), .eq(weq576));
    equaln #(12) e577(.a(buffered_input), .b(12'b001001000001), .eq(weq577));
    equaln #(12) e578(.a(buffered_input), .b(12'b001001000010), .eq(weq578));
    equaln #(12) e579(.a(buffered_input), .b(12'b001001000011), .eq(weq579));
    equaln #(12) e580(.a(buffered_input), .b(12'b001001000100), .eq(weq580));
    equaln #(12) e581(.a(buffered_input), .b(12'b001001000101), .eq(weq581));
    equaln #(12) e582(.a(buffered_input), .b(12'b001001000110), .eq(weq582));
    equaln #(12) e583(.a(buffered_input), .b(12'b001001000111), .eq(weq583));
    equaln #(12) e584(.a(buffered_input), .b(12'b001001001000), .eq(weq584));
    equaln #(12) e585(.a(buffered_input), .b(12'b001001001001), .eq(weq585));
    equaln #(12) e586(.a(buffered_input), .b(12'b001001001010), .eq(weq586));
    equaln #(12) e587(.a(buffered_input), .b(12'b001001001011), .eq(weq587));
    equaln #(12) e588(.a(buffered_input), .b(12'b001001001100), .eq(weq588));
    equaln #(12) e589(.a(buffered_input), .b(12'b001001001101), .eq(weq589));
    equaln #(12) e590(.a(buffered_input), .b(12'b001001001110), .eq(weq590));
    equaln #(12) e591(.a(buffered_input), .b(12'b001001001111), .eq(weq591));
    equaln #(12) e592(.a(buffered_input), .b(12'b001001010000), .eq(weq592));
    equaln #(12) e593(.a(buffered_input), .b(12'b001001010001), .eq(weq593));
    equaln #(12) e594(.a(buffered_input), .b(12'b001001010010), .eq(weq594));
    equaln #(12) e595(.a(buffered_input), .b(12'b001001010011), .eq(weq595));
    equaln #(12) e596(.a(buffered_input), .b(12'b001001010100), .eq(weq596));
    equaln #(12) e597(.a(buffered_input), .b(12'b001001010101), .eq(weq597));
    equaln #(12) e598(.a(buffered_input), .b(12'b001001010110), .eq(weq598));
    equaln #(12) e599(.a(buffered_input), .b(12'b001001010111), .eq(weq599));
    equaln #(12) e600(.a(buffered_input), .b(12'b001001011000), .eq(weq600));
    equaln #(12) e601(.a(buffered_input), .b(12'b001001011001), .eq(weq601));
    equaln #(12) e602(.a(buffered_input), .b(12'b001001011010), .eq(weq602));
    equaln #(12) e603(.a(buffered_input), .b(12'b001001011011), .eq(weq603));
    equaln #(12) e604(.a(buffered_input), .b(12'b001001011100), .eq(weq604));
    equaln #(12) e605(.a(buffered_input), .b(12'b001001011101), .eq(weq605));
    equaln #(12) e606(.a(buffered_input), .b(12'b001001011110), .eq(weq606));
    equaln #(12) e607(.a(buffered_input), .b(12'b001001011111), .eq(weq607));
    equaln #(12) e608(.a(buffered_input), .b(12'b001001100000), .eq(weq608));
    equaln #(12) e609(.a(buffered_input), .b(12'b001001100001), .eq(weq609));
    equaln #(12) e610(.a(buffered_input), .b(12'b001001100010), .eq(weq610));
    equaln #(12) e611(.a(buffered_input), .b(12'b001001100011), .eq(weq611));
    equaln #(12) e612(.a(buffered_input), .b(12'b001001100100), .eq(weq612));
    equaln #(12) e613(.a(buffered_input), .b(12'b001001100101), .eq(weq613));
    equaln #(12) e614(.a(buffered_input), .b(12'b001001100110), .eq(weq614));
    equaln #(12) e615(.a(buffered_input), .b(12'b001001100111), .eq(weq615));
    equaln #(12) e616(.a(buffered_input), .b(12'b001001101000), .eq(weq616));
    equaln #(12) e617(.a(buffered_input), .b(12'b001001101001), .eq(weq617));
    equaln #(12) e618(.a(buffered_input), .b(12'b001001101010), .eq(weq618));
    equaln #(12) e619(.a(buffered_input), .b(12'b001001101011), .eq(weq619));
    equaln #(12) e620(.a(buffered_input), .b(12'b001001101100), .eq(weq620));
    equaln #(12) e621(.a(buffered_input), .b(12'b001001101101), .eq(weq621));
    equaln #(12) e622(.a(buffered_input), .b(12'b001001101110), .eq(weq622));
    equaln #(12) e623(.a(buffered_input), .b(12'b001001101111), .eq(weq623));
    equaln #(12) e624(.a(buffered_input), .b(12'b001001110000), .eq(weq624));
    equaln #(12) e625(.a(buffered_input), .b(12'b001001110001), .eq(weq625));
    equaln #(12) e626(.a(buffered_input), .b(12'b001001110010), .eq(weq626));
    equaln #(12) e627(.a(buffered_input), .b(12'b001001110011), .eq(weq627));
    equaln #(12) e628(.a(buffered_input), .b(12'b001001110100), .eq(weq628));
    equaln #(12) e629(.a(buffered_input), .b(12'b001001110101), .eq(weq629));
    equaln #(12) e630(.a(buffered_input), .b(12'b001001110110), .eq(weq630));
    equaln #(12) e631(.a(buffered_input), .b(12'b001001110111), .eq(weq631));
    equaln #(12) e632(.a(buffered_input), .b(12'b001001111000), .eq(weq632));
    equaln #(12) e633(.a(buffered_input), .b(12'b001001111001), .eq(weq633));
    equaln #(12) e634(.a(buffered_input), .b(12'b001001111010), .eq(weq634));
    equaln #(12) e635(.a(buffered_input), .b(12'b001001111011), .eq(weq635));
    equaln #(12) e636(.a(buffered_input), .b(12'b001001111100), .eq(weq636));
    equaln #(12) e637(.a(buffered_input), .b(12'b001001111101), .eq(weq637));
    equaln #(12) e638(.a(buffered_input), .b(12'b001001111110), .eq(weq638));
    equaln #(12) e639(.a(buffered_input), .b(12'b001001111111), .eq(weq639));
    equaln #(12) e640(.a(buffered_input), .b(12'b001010000000), .eq(weq640));
    equaln #(12) e641(.a(buffered_input), .b(12'b001010000001), .eq(weq641));
    equaln #(12) e642(.a(buffered_input), .b(12'b001010000010), .eq(weq642));
    equaln #(12) e643(.a(buffered_input), .b(12'b001010000011), .eq(weq643));
    equaln #(12) e644(.a(buffered_input), .b(12'b001010000100), .eq(weq644));
    equaln #(12) e645(.a(buffered_input), .b(12'b001010000101), .eq(weq645));
    equaln #(12) e646(.a(buffered_input), .b(12'b001010000110), .eq(weq646));
    equaln #(12) e647(.a(buffered_input), .b(12'b001010000111), .eq(weq647));
    equaln #(12) e648(.a(buffered_input), .b(12'b001010001000), .eq(weq648));
    equaln #(12) e649(.a(buffered_input), .b(12'b001010001001), .eq(weq649));
    equaln #(12) e650(.a(buffered_input), .b(12'b001010001010), .eq(weq650));
    equaln #(12) e651(.a(buffered_input), .b(12'b001010001011), .eq(weq651));
    equaln #(12) e652(.a(buffered_input), .b(12'b001010001100), .eq(weq652));
    equaln #(12) e653(.a(buffered_input), .b(12'b001010001101), .eq(weq653));
    equaln #(12) e654(.a(buffered_input), .b(12'b001010001110), .eq(weq654));
    equaln #(12) e655(.a(buffered_input), .b(12'b001010001111), .eq(weq655));
    equaln #(12) e656(.a(buffered_input), .b(12'b001010010000), .eq(weq656));
    equaln #(12) e657(.a(buffered_input), .b(12'b001010010001), .eq(weq657));
    equaln #(12) e658(.a(buffered_input), .b(12'b001010010010), .eq(weq658));
    equaln #(12) e659(.a(buffered_input), .b(12'b001010010011), .eq(weq659));
    equaln #(12) e660(.a(buffered_input), .b(12'b001010010100), .eq(weq660));
    equaln #(12) e661(.a(buffered_input), .b(12'b001010010101), .eq(weq661));
    equaln #(12) e662(.a(buffered_input), .b(12'b001010010110), .eq(weq662));
    equaln #(12) e663(.a(buffered_input), .b(12'b001010010111), .eq(weq663));
    equaln #(12) e664(.a(buffered_input), .b(12'b001010011000), .eq(weq664));
    equaln #(12) e665(.a(buffered_input), .b(12'b001010011001), .eq(weq665));
    equaln #(12) e666(.a(buffered_input), .b(12'b001010011010), .eq(weq666));
    equaln #(12) e667(.a(buffered_input), .b(12'b001010011011), .eq(weq667));
    equaln #(12) e668(.a(buffered_input), .b(12'b001010011100), .eq(weq668));
    equaln #(12) e669(.a(buffered_input), .b(12'b001010011101), .eq(weq669));
    equaln #(12) e670(.a(buffered_input), .b(12'b001010011110), .eq(weq670));
    equaln #(12) e671(.a(buffered_input), .b(12'b001010011111), .eq(weq671));
    equaln #(12) e672(.a(buffered_input), .b(12'b001010100000), .eq(weq672));
    equaln #(12) e673(.a(buffered_input), .b(12'b001010100001), .eq(weq673));
    equaln #(12) e674(.a(buffered_input), .b(12'b001010100010), .eq(weq674));
    equaln #(12) e675(.a(buffered_input), .b(12'b001010100011), .eq(weq675));
    equaln #(12) e676(.a(buffered_input), .b(12'b001010100100), .eq(weq676));
    equaln #(12) e677(.a(buffered_input), .b(12'b001010100101), .eq(weq677));
    equaln #(12) e678(.a(buffered_input), .b(12'b001010100110), .eq(weq678));
    equaln #(12) e679(.a(buffered_input), .b(12'b001010100111), .eq(weq679));
    equaln #(12) e680(.a(buffered_input), .b(12'b001010101000), .eq(weq680));
    equaln #(12) e681(.a(buffered_input), .b(12'b001010101001), .eq(weq681));
    equaln #(12) e682(.a(buffered_input), .b(12'b001010101010), .eq(weq682));
    equaln #(12) e683(.a(buffered_input), .b(12'b001010101011), .eq(weq683));
    equaln #(12) e684(.a(buffered_input), .b(12'b001010101100), .eq(weq684));
    equaln #(12) e685(.a(buffered_input), .b(12'b001010101101), .eq(weq685));
    equaln #(12) e686(.a(buffered_input), .b(12'b001010101110), .eq(weq686));
    equaln #(12) e687(.a(buffered_input), .b(12'b001010101111), .eq(weq687));
    equaln #(12) e688(.a(buffered_input), .b(12'b001010110000), .eq(weq688));
    equaln #(12) e689(.a(buffered_input), .b(12'b001010110001), .eq(weq689));
    equaln #(12) e690(.a(buffered_input), .b(12'b001010110010), .eq(weq690));
    equaln #(12) e691(.a(buffered_input), .b(12'b001010110011), .eq(weq691));
    equaln #(12) e692(.a(buffered_input), .b(12'b001010110100), .eq(weq692));
    equaln #(12) e693(.a(buffered_input), .b(12'b001010110101), .eq(weq693));
    equaln #(12) e694(.a(buffered_input), .b(12'b001010110110), .eq(weq694));
    equaln #(12) e695(.a(buffered_input), .b(12'b001010110111), .eq(weq695));
    equaln #(12) e696(.a(buffered_input), .b(12'b001010111000), .eq(weq696));
    equaln #(12) e697(.a(buffered_input), .b(12'b001010111001), .eq(weq697));
    equaln #(12) e698(.a(buffered_input), .b(12'b001010111010), .eq(weq698));
    equaln #(12) e699(.a(buffered_input), .b(12'b001010111011), .eq(weq699));
    equaln #(12) e700(.a(buffered_input), .b(12'b001010111100), .eq(weq700));
    equaln #(12) e701(.a(buffered_input), .b(12'b001010111101), .eq(weq701));
    equaln #(12) e702(.a(buffered_input), .b(12'b001010111110), .eq(weq702));
    equaln #(12) e703(.a(buffered_input), .b(12'b001010111111), .eq(weq703));
    equaln #(12) e704(.a(buffered_input), .b(12'b001011000000), .eq(weq704));
    equaln #(12) e705(.a(buffered_input), .b(12'b001011000001), .eq(weq705));
    equaln #(12) e706(.a(buffered_input), .b(12'b001011000010), .eq(weq706));
    equaln #(12) e707(.a(buffered_input), .b(12'b001011000011), .eq(weq707));
    equaln #(12) e708(.a(buffered_input), .b(12'b001011000100), .eq(weq708));
    equaln #(12) e709(.a(buffered_input), .b(12'b001011000101), .eq(weq709));
    equaln #(12) e710(.a(buffered_input), .b(12'b001011000110), .eq(weq710));
    equaln #(12) e711(.a(buffered_input), .b(12'b001011000111), .eq(weq711));
    equaln #(12) e712(.a(buffered_input), .b(12'b001011001000), .eq(weq712));
    equaln #(12) e713(.a(buffered_input), .b(12'b001011001001), .eq(weq713));
    equaln #(12) e714(.a(buffered_input), .b(12'b001011001010), .eq(weq714));
    equaln #(12) e715(.a(buffered_input), .b(12'b001011001011), .eq(weq715));
    equaln #(12) e716(.a(buffered_input), .b(12'b001011001100), .eq(weq716));
    equaln #(12) e717(.a(buffered_input), .b(12'b001011001101), .eq(weq717));
    equaln #(12) e718(.a(buffered_input), .b(12'b001011001110), .eq(weq718));
    equaln #(12) e719(.a(buffered_input), .b(12'b001011001111), .eq(weq719));
    equaln #(12) e720(.a(buffered_input), .b(12'b001011010000), .eq(weq720));
    equaln #(12) e721(.a(buffered_input), .b(12'b001011010001), .eq(weq721));
    equaln #(12) e722(.a(buffered_input), .b(12'b001011010010), .eq(weq722));
    equaln #(12) e723(.a(buffered_input), .b(12'b001011010011), .eq(weq723));
    equaln #(12) e724(.a(buffered_input), .b(12'b001011010100), .eq(weq724));
    equaln #(12) e725(.a(buffered_input), .b(12'b001011010101), .eq(weq725));
    equaln #(12) e726(.a(buffered_input), .b(12'b001011010110), .eq(weq726));
    equaln #(12) e727(.a(buffered_input), .b(12'b001011010111), .eq(weq727));
    equaln #(12) e728(.a(buffered_input), .b(12'b001011011000), .eq(weq728));
    equaln #(12) e729(.a(buffered_input), .b(12'b001011011001), .eq(weq729));
    equaln #(12) e730(.a(buffered_input), .b(12'b001011011010), .eq(weq730));
    equaln #(12) e731(.a(buffered_input), .b(12'b001011011011), .eq(weq731));
    equaln #(12) e732(.a(buffered_input), .b(12'b001011011100), .eq(weq732));
    equaln #(12) e733(.a(buffered_input), .b(12'b001011011101), .eq(weq733));
    equaln #(12) e734(.a(buffered_input), .b(12'b001011011110), .eq(weq734));
    equaln #(12) e735(.a(buffered_input), .b(12'b001011011111), .eq(weq735));
    equaln #(12) e736(.a(buffered_input), .b(12'b001011100000), .eq(weq736));
    equaln #(12) e737(.a(buffered_input), .b(12'b001011100001), .eq(weq737));
    equaln #(12) e738(.a(buffered_input), .b(12'b001011100010), .eq(weq738));
    equaln #(12) e739(.a(buffered_input), .b(12'b001011100011), .eq(weq739));
    equaln #(12) e740(.a(buffered_input), .b(12'b001011100100), .eq(weq740));
    equaln #(12) e741(.a(buffered_input), .b(12'b001011100101), .eq(weq741));
    equaln #(12) e742(.a(buffered_input), .b(12'b001011100110), .eq(weq742));
    equaln #(12) e743(.a(buffered_input), .b(12'b001011100111), .eq(weq743));
    equaln #(12) e744(.a(buffered_input), .b(12'b001011101000), .eq(weq744));
    equaln #(12) e745(.a(buffered_input), .b(12'b001011101001), .eq(weq745));
    equaln #(12) e746(.a(buffered_input), .b(12'b001011101010), .eq(weq746));
    equaln #(12) e747(.a(buffered_input), .b(12'b001011101011), .eq(weq747));
    equaln #(12) e748(.a(buffered_input), .b(12'b001011101100), .eq(weq748));
    equaln #(12) e749(.a(buffered_input), .b(12'b001011101101), .eq(weq749));
    equaln #(12) e750(.a(buffered_input), .b(12'b001011101110), .eq(weq750));
    equaln #(12) e751(.a(buffered_input), .b(12'b001011101111), .eq(weq751));
    equaln #(12) e752(.a(buffered_input), .b(12'b001011110000), .eq(weq752));
    equaln #(12) e753(.a(buffered_input), .b(12'b001011110001), .eq(weq753));
    equaln #(12) e754(.a(buffered_input), .b(12'b001011110010), .eq(weq754));
    equaln #(12) e755(.a(buffered_input), .b(12'b001011110011), .eq(weq755));
    equaln #(12) e756(.a(buffered_input), .b(12'b001011110100), .eq(weq756));
    equaln #(12) e757(.a(buffered_input), .b(12'b001011110101), .eq(weq757));
    equaln #(12) e758(.a(buffered_input), .b(12'b001011110110), .eq(weq758));
    equaln #(12) e759(.a(buffered_input), .b(12'b001011110111), .eq(weq759));
    equaln #(12) e760(.a(buffered_input), .b(12'b001011111000), .eq(weq760));
    equaln #(12) e761(.a(buffered_input), .b(12'b001011111001), .eq(weq761));
    equaln #(12) e762(.a(buffered_input), .b(12'b001011111010), .eq(weq762));
    equaln #(12) e763(.a(buffered_input), .b(12'b001011111011), .eq(weq763));
    equaln #(12) e764(.a(buffered_input), .b(12'b001011111100), .eq(weq764));
    equaln #(12) e765(.a(buffered_input), .b(12'b001011111101), .eq(weq765));
    equaln #(12) e766(.a(buffered_input), .b(12'b001011111110), .eq(weq766));
    equaln #(12) e767(.a(buffered_input), .b(12'b001011111111), .eq(weq767));
    equaln #(12) e768(.a(buffered_input), .b(12'b001100000000), .eq(weq768));
    equaln #(12) e769(.a(buffered_input), .b(12'b001100000001), .eq(weq769));
    equaln #(12) e770(.a(buffered_input), .b(12'b001100000010), .eq(weq770));
    equaln #(12) e771(.a(buffered_input), .b(12'b001100000011), .eq(weq771));
    equaln #(12) e772(.a(buffered_input), .b(12'b001100000100), .eq(weq772));
    equaln #(12) e773(.a(buffered_input), .b(12'b001100000101), .eq(weq773));
    equaln #(12) e774(.a(buffered_input), .b(12'b001100000110), .eq(weq774));
    equaln #(12) e775(.a(buffered_input), .b(12'b001100000111), .eq(weq775));
    equaln #(12) e776(.a(buffered_input), .b(12'b001100001000), .eq(weq776));
    equaln #(12) e777(.a(buffered_input), .b(12'b001100001001), .eq(weq777));
    equaln #(12) e778(.a(buffered_input), .b(12'b001100001010), .eq(weq778));
    equaln #(12) e779(.a(buffered_input), .b(12'b001100001011), .eq(weq779));
    equaln #(12) e780(.a(buffered_input), .b(12'b001100001100), .eq(weq780));
    equaln #(12) e781(.a(buffered_input), .b(12'b001100001101), .eq(weq781));
    equaln #(12) e782(.a(buffered_input), .b(12'b001100001110), .eq(weq782));
    equaln #(12) e783(.a(buffered_input), .b(12'b001100001111), .eq(weq783));
    equaln #(12) e784(.a(buffered_input), .b(12'b001100010000), .eq(weq784));
    equaln #(12) e785(.a(buffered_input), .b(12'b001100010001), .eq(weq785));
    equaln #(12) e786(.a(buffered_input), .b(12'b001100010010), .eq(weq786));
    equaln #(12) e787(.a(buffered_input), .b(12'b001100010011), .eq(weq787));
    equaln #(12) e788(.a(buffered_input), .b(12'b001100010100), .eq(weq788));
    equaln #(12) e789(.a(buffered_input), .b(12'b001100010101), .eq(weq789));
    equaln #(12) e790(.a(buffered_input), .b(12'b001100010110), .eq(weq790));
    equaln #(12) e791(.a(buffered_input), .b(12'b001100010111), .eq(weq791));
    equaln #(12) e792(.a(buffered_input), .b(12'b001100011000), .eq(weq792));
    equaln #(12) e793(.a(buffered_input), .b(12'b001100011001), .eq(weq793));
    equaln #(12) e794(.a(buffered_input), .b(12'b001100011010), .eq(weq794));
    equaln #(12) e795(.a(buffered_input), .b(12'b001100011011), .eq(weq795));
    equaln #(12) e796(.a(buffered_input), .b(12'b001100011100), .eq(weq796));
    equaln #(12) e797(.a(buffered_input), .b(12'b001100011101), .eq(weq797));
    equaln #(12) e798(.a(buffered_input), .b(12'b001100011110), .eq(weq798));
    equaln #(12) e799(.a(buffered_input), .b(12'b001100011111), .eq(weq799));
    equaln #(12) e800(.a(buffered_input), .b(12'b001100100000), .eq(weq800));
    equaln #(12) e801(.a(buffered_input), .b(12'b001100100001), .eq(weq801));
    equaln #(12) e802(.a(buffered_input), .b(12'b001100100010), .eq(weq802));
    equaln #(12) e803(.a(buffered_input), .b(12'b001100100011), .eq(weq803));
    equaln #(12) e804(.a(buffered_input), .b(12'b001100100100), .eq(weq804));
    equaln #(12) e805(.a(buffered_input), .b(12'b001100100101), .eq(weq805));
    equaln #(12) e806(.a(buffered_input), .b(12'b001100100110), .eq(weq806));
    equaln #(12) e807(.a(buffered_input), .b(12'b001100100111), .eq(weq807));
    equaln #(12) e808(.a(buffered_input), .b(12'b001100101000), .eq(weq808));
    equaln #(12) e809(.a(buffered_input), .b(12'b001100101001), .eq(weq809));
    equaln #(12) e810(.a(buffered_input), .b(12'b001100101010), .eq(weq810));
    equaln #(12) e811(.a(buffered_input), .b(12'b001100101011), .eq(weq811));
    equaln #(12) e812(.a(buffered_input), .b(12'b001100101100), .eq(weq812));
    equaln #(12) e813(.a(buffered_input), .b(12'b001100101101), .eq(weq813));
    equaln #(12) e814(.a(buffered_input), .b(12'b001100101110), .eq(weq814));
    equaln #(12) e815(.a(buffered_input), .b(12'b001100101111), .eq(weq815));
    equaln #(12) e816(.a(buffered_input), .b(12'b001100110000), .eq(weq816));
    equaln #(12) e817(.a(buffered_input), .b(12'b001100110001), .eq(weq817));
    equaln #(12) e818(.a(buffered_input), .b(12'b001100110010), .eq(weq818));
    equaln #(12) e819(.a(buffered_input), .b(12'b001100110011), .eq(weq819));
    equaln #(12) e820(.a(buffered_input), .b(12'b001100110100), .eq(weq820));
    equaln #(12) e821(.a(buffered_input), .b(12'b001100110101), .eq(weq821));
    equaln #(12) e822(.a(buffered_input), .b(12'b001100110110), .eq(weq822));
    equaln #(12) e823(.a(buffered_input), .b(12'b001100110111), .eq(weq823));
    equaln #(12) e824(.a(buffered_input), .b(12'b001100111000), .eq(weq824));
    equaln #(12) e825(.a(buffered_input), .b(12'b001100111001), .eq(weq825));
    equaln #(12) e826(.a(buffered_input), .b(12'b001100111010), .eq(weq826));
    equaln #(12) e827(.a(buffered_input), .b(12'b001100111011), .eq(weq827));
    equaln #(12) e828(.a(buffered_input), .b(12'b001100111100), .eq(weq828));
    equaln #(12) e829(.a(buffered_input), .b(12'b001100111101), .eq(weq829));
    equaln #(12) e830(.a(buffered_input), .b(12'b001100111110), .eq(weq830));
    equaln #(12) e831(.a(buffered_input), .b(12'b001100111111), .eq(weq831));
    equaln #(12) e832(.a(buffered_input), .b(12'b001101000000), .eq(weq832));
    equaln #(12) e833(.a(buffered_input), .b(12'b001101000001), .eq(weq833));
    equaln #(12) e834(.a(buffered_input), .b(12'b001101000010), .eq(weq834));
    equaln #(12) e835(.a(buffered_input), .b(12'b001101000011), .eq(weq835));
    equaln #(12) e836(.a(buffered_input), .b(12'b001101000100), .eq(weq836));
    equaln #(12) e837(.a(buffered_input), .b(12'b001101000101), .eq(weq837));
    equaln #(12) e838(.a(buffered_input), .b(12'b001101000110), .eq(weq838));
    equaln #(12) e839(.a(buffered_input), .b(12'b001101000111), .eq(weq839));
    equaln #(12) e840(.a(buffered_input), .b(12'b001101001000), .eq(weq840));
    equaln #(12) e841(.a(buffered_input), .b(12'b001101001001), .eq(weq841));
    equaln #(12) e842(.a(buffered_input), .b(12'b001101001010), .eq(weq842));
    equaln #(12) e843(.a(buffered_input), .b(12'b001101001011), .eq(weq843));
    equaln #(12) e844(.a(buffered_input), .b(12'b001101001100), .eq(weq844));
    equaln #(12) e845(.a(buffered_input), .b(12'b001101001101), .eq(weq845));
    equaln #(12) e846(.a(buffered_input), .b(12'b001101001110), .eq(weq846));
    equaln #(12) e847(.a(buffered_input), .b(12'b001101001111), .eq(weq847));
    equaln #(12) e848(.a(buffered_input), .b(12'b001101010000), .eq(weq848));
    equaln #(12) e849(.a(buffered_input), .b(12'b001101010001), .eq(weq849));
    equaln #(12) e850(.a(buffered_input), .b(12'b001101010010), .eq(weq850));
    equaln #(12) e851(.a(buffered_input), .b(12'b001101010011), .eq(weq851));
    equaln #(12) e852(.a(buffered_input), .b(12'b001101010100), .eq(weq852));
    equaln #(12) e853(.a(buffered_input), .b(12'b001101010101), .eq(weq853));
    equaln #(12) e854(.a(buffered_input), .b(12'b001101010110), .eq(weq854));
    equaln #(12) e855(.a(buffered_input), .b(12'b001101010111), .eq(weq855));
    equaln #(12) e856(.a(buffered_input), .b(12'b001101011000), .eq(weq856));
    equaln #(12) e857(.a(buffered_input), .b(12'b001101011001), .eq(weq857));
    equaln #(12) e858(.a(buffered_input), .b(12'b001101011010), .eq(weq858));
    equaln #(12) e859(.a(buffered_input), .b(12'b001101011011), .eq(weq859));
    equaln #(12) e860(.a(buffered_input), .b(12'b001101011100), .eq(weq860));
    equaln #(12) e861(.a(buffered_input), .b(12'b001101011101), .eq(weq861));
    equaln #(12) e862(.a(buffered_input), .b(12'b001101011110), .eq(weq862));
    equaln #(12) e863(.a(buffered_input), .b(12'b001101011111), .eq(weq863));
    equaln #(12) e864(.a(buffered_input), .b(12'b001101100000), .eq(weq864));
    equaln #(12) e865(.a(buffered_input), .b(12'b001101100001), .eq(weq865));
    equaln #(12) e866(.a(buffered_input), .b(12'b001101100010), .eq(weq866));
    equaln #(12) e867(.a(buffered_input), .b(12'b001101100011), .eq(weq867));
    equaln #(12) e868(.a(buffered_input), .b(12'b001101100100), .eq(weq868));
    equaln #(12) e869(.a(buffered_input), .b(12'b001101100101), .eq(weq869));
    equaln #(12) e870(.a(buffered_input), .b(12'b001101100110), .eq(weq870));
    equaln #(12) e871(.a(buffered_input), .b(12'b001101100111), .eq(weq871));
    equaln #(12) e872(.a(buffered_input), .b(12'b001101101000), .eq(weq872));
    equaln #(12) e873(.a(buffered_input), .b(12'b001101101001), .eq(weq873));
    equaln #(12) e874(.a(buffered_input), .b(12'b001101101010), .eq(weq874));
    equaln #(12) e875(.a(buffered_input), .b(12'b001101101011), .eq(weq875));
    equaln #(12) e876(.a(buffered_input), .b(12'b001101101100), .eq(weq876));
    equaln #(12) e877(.a(buffered_input), .b(12'b001101101101), .eq(weq877));
    equaln #(12) e878(.a(buffered_input), .b(12'b001101101110), .eq(weq878));
    equaln #(12) e879(.a(buffered_input), .b(12'b001101101111), .eq(weq879));
    equaln #(12) e880(.a(buffered_input), .b(12'b001101110000), .eq(weq880));
    equaln #(12) e881(.a(buffered_input), .b(12'b001101110001), .eq(weq881));
    equaln #(12) e882(.a(buffered_input), .b(12'b001101110010), .eq(weq882));
    equaln #(12) e883(.a(buffered_input), .b(12'b001101110011), .eq(weq883));
    equaln #(12) e884(.a(buffered_input), .b(12'b001101110100), .eq(weq884));
    equaln #(12) e885(.a(buffered_input), .b(12'b001101110101), .eq(weq885));
    equaln #(12) e886(.a(buffered_input), .b(12'b001101110110), .eq(weq886));
    equaln #(12) e887(.a(buffered_input), .b(12'b001101110111), .eq(weq887));
    equaln #(12) e888(.a(buffered_input), .b(12'b001101111000), .eq(weq888));
    equaln #(12) e889(.a(buffered_input), .b(12'b001101111001), .eq(weq889));
    equaln #(12) e890(.a(buffered_input), .b(12'b001101111010), .eq(weq890));
    equaln #(12) e891(.a(buffered_input), .b(12'b001101111011), .eq(weq891));
    equaln #(12) e892(.a(buffered_input), .b(12'b001101111100), .eq(weq892));
    equaln #(12) e893(.a(buffered_input), .b(12'b001101111101), .eq(weq893));
    equaln #(12) e894(.a(buffered_input), .b(12'b001101111110), .eq(weq894));
    equaln #(12) e895(.a(buffered_input), .b(12'b001101111111), .eq(weq895));
    equaln #(12) e896(.a(buffered_input), .b(12'b001110000000), .eq(weq896));
    equaln #(12) e897(.a(buffered_input), .b(12'b001110000001), .eq(weq897));
    equaln #(12) e898(.a(buffered_input), .b(12'b001110000010), .eq(weq898));
    equaln #(12) e899(.a(buffered_input), .b(12'b001110000011), .eq(weq899));
    equaln #(12) e900(.a(buffered_input), .b(12'b001110000100), .eq(weq900));
    equaln #(12) e901(.a(buffered_input), .b(12'b001110000101), .eq(weq901));
    equaln #(12) e902(.a(buffered_input), .b(12'b001110000110), .eq(weq902));
    equaln #(12) e903(.a(buffered_input), .b(12'b001110000111), .eq(weq903));
    equaln #(12) e904(.a(buffered_input), .b(12'b001110001000), .eq(weq904));
    equaln #(12) e905(.a(buffered_input), .b(12'b001110001001), .eq(weq905));
    equaln #(12) e906(.a(buffered_input), .b(12'b001110001010), .eq(weq906));
    equaln #(12) e907(.a(buffered_input), .b(12'b001110001011), .eq(weq907));
    equaln #(12) e908(.a(buffered_input), .b(12'b001110001100), .eq(weq908));
    equaln #(12) e909(.a(buffered_input), .b(12'b001110001101), .eq(weq909));
    equaln #(12) e910(.a(buffered_input), .b(12'b001110001110), .eq(weq910));
    equaln #(12) e911(.a(buffered_input), .b(12'b001110001111), .eq(weq911));
    equaln #(12) e912(.a(buffered_input), .b(12'b001110010000), .eq(weq912));
    equaln #(12) e913(.a(buffered_input), .b(12'b001110010001), .eq(weq913));
    equaln #(12) e914(.a(buffered_input), .b(12'b001110010010), .eq(weq914));
    equaln #(12) e915(.a(buffered_input), .b(12'b001110010011), .eq(weq915));
    equaln #(12) e916(.a(buffered_input), .b(12'b001110010100), .eq(weq916));
    equaln #(12) e917(.a(buffered_input), .b(12'b001110010101), .eq(weq917));
    equaln #(12) e918(.a(buffered_input), .b(12'b001110010110), .eq(weq918));
    equaln #(12) e919(.a(buffered_input), .b(12'b001110010111), .eq(weq919));
    equaln #(12) e920(.a(buffered_input), .b(12'b001110011000), .eq(weq920));
    equaln #(12) e921(.a(buffered_input), .b(12'b001110011001), .eq(weq921));
    equaln #(12) e922(.a(buffered_input), .b(12'b001110011010), .eq(weq922));
    equaln #(12) e923(.a(buffered_input), .b(12'b001110011011), .eq(weq923));
    equaln #(12) e924(.a(buffered_input), .b(12'b001110011100), .eq(weq924));
    equaln #(12) e925(.a(buffered_input), .b(12'b001110011101), .eq(weq925));
    equaln #(12) e926(.a(buffered_input), .b(12'b001110011110), .eq(weq926));
    equaln #(12) e927(.a(buffered_input), .b(12'b001110011111), .eq(weq927));
    equaln #(12) e928(.a(buffered_input), .b(12'b001110100000), .eq(weq928));
    equaln #(12) e929(.a(buffered_input), .b(12'b001110100001), .eq(weq929));
    equaln #(12) e930(.a(buffered_input), .b(12'b001110100010), .eq(weq930));
    equaln #(12) e931(.a(buffered_input), .b(12'b001110100011), .eq(weq931));
    equaln #(12) e932(.a(buffered_input), .b(12'b001110100100), .eq(weq932));
    equaln #(12) e933(.a(buffered_input), .b(12'b001110100101), .eq(weq933));
    equaln #(12) e934(.a(buffered_input), .b(12'b001110100110), .eq(weq934));
    equaln #(12) e935(.a(buffered_input), .b(12'b001110100111), .eq(weq935));
    equaln #(12) e936(.a(buffered_input), .b(12'b001110101000), .eq(weq936));
    equaln #(12) e937(.a(buffered_input), .b(12'b001110101001), .eq(weq937));
    equaln #(12) e938(.a(buffered_input), .b(12'b001110101010), .eq(weq938));
    equaln #(12) e939(.a(buffered_input), .b(12'b001110101011), .eq(weq939));
    equaln #(12) e940(.a(buffered_input), .b(12'b001110101100), .eq(weq940));
    equaln #(12) e941(.a(buffered_input), .b(12'b001110101101), .eq(weq941));
    equaln #(12) e942(.a(buffered_input), .b(12'b001110101110), .eq(weq942));
    equaln #(12) e943(.a(buffered_input), .b(12'b001110101111), .eq(weq943));
    equaln #(12) e944(.a(buffered_input), .b(12'b001110110000), .eq(weq944));
    equaln #(12) e945(.a(buffered_input), .b(12'b001110110001), .eq(weq945));
    equaln #(12) e946(.a(buffered_input), .b(12'b001110110010), .eq(weq946));
    equaln #(12) e947(.a(buffered_input), .b(12'b001110110011), .eq(weq947));
    equaln #(12) e948(.a(buffered_input), .b(12'b001110110100), .eq(weq948));
    equaln #(12) e949(.a(buffered_input), .b(12'b001110110101), .eq(weq949));
    equaln #(12) e950(.a(buffered_input), .b(12'b001110110110), .eq(weq950));
    equaln #(12) e951(.a(buffered_input), .b(12'b001110110111), .eq(weq951));
    equaln #(12) e952(.a(buffered_input), .b(12'b001110111000), .eq(weq952));
    equaln #(12) e953(.a(buffered_input), .b(12'b001110111001), .eq(weq953));
    equaln #(12) e954(.a(buffered_input), .b(12'b001110111010), .eq(weq954));
    equaln #(12) e955(.a(buffered_input), .b(12'b001110111011), .eq(weq955));
    equaln #(12) e956(.a(buffered_input), .b(12'b001110111100), .eq(weq956));
    equaln #(12) e957(.a(buffered_input), .b(12'b001110111101), .eq(weq957));
    equaln #(12) e958(.a(buffered_input), .b(12'b001110111110), .eq(weq958));
    equaln #(12) e959(.a(buffered_input), .b(12'b001110111111), .eq(weq959));
    equaln #(12) e960(.a(buffered_input), .b(12'b001111000000), .eq(weq960));
    equaln #(12) e961(.a(buffered_input), .b(12'b001111000001), .eq(weq961));
    equaln #(12) e962(.a(buffered_input), .b(12'b001111000010), .eq(weq962));
    equaln #(12) e963(.a(buffered_input), .b(12'b001111000011), .eq(weq963));
    equaln #(12) e964(.a(buffered_input), .b(12'b001111000100), .eq(weq964));
    equaln #(12) e965(.a(buffered_input), .b(12'b001111000101), .eq(weq965));
    equaln #(12) e966(.a(buffered_input), .b(12'b001111000110), .eq(weq966));
    equaln #(12) e967(.a(buffered_input), .b(12'b001111000111), .eq(weq967));
    equaln #(12) e968(.a(buffered_input), .b(12'b001111001000), .eq(weq968));
    equaln #(12) e969(.a(buffered_input), .b(12'b001111001001), .eq(weq969));
    equaln #(12) e970(.a(buffered_input), .b(12'b001111001010), .eq(weq970));
    equaln #(12) e971(.a(buffered_input), .b(12'b001111001011), .eq(weq971));
    equaln #(12) e972(.a(buffered_input), .b(12'b001111001100), .eq(weq972));
    equaln #(12) e973(.a(buffered_input), .b(12'b001111001101), .eq(weq973));
    equaln #(12) e974(.a(buffered_input), .b(12'b001111001110), .eq(weq974));
    equaln #(12) e975(.a(buffered_input), .b(12'b001111001111), .eq(weq975));
    equaln #(12) e976(.a(buffered_input), .b(12'b001111010000), .eq(weq976));
    equaln #(12) e977(.a(buffered_input), .b(12'b001111010001), .eq(weq977));
    equaln #(12) e978(.a(buffered_input), .b(12'b001111010010), .eq(weq978));
    equaln #(12) e979(.a(buffered_input), .b(12'b001111010011), .eq(weq979));
    equaln #(12) e980(.a(buffered_input), .b(12'b001111010100), .eq(weq980));
    equaln #(12) e981(.a(buffered_input), .b(12'b001111010101), .eq(weq981));
    equaln #(12) e982(.a(buffered_input), .b(12'b001111010110), .eq(weq982));
    equaln #(12) e983(.a(buffered_input), .b(12'b001111010111), .eq(weq983));
    equaln #(12) e984(.a(buffered_input), .b(12'b001111011000), .eq(weq984));
    equaln #(12) e985(.a(buffered_input), .b(12'b001111011001), .eq(weq985));
    equaln #(12) e986(.a(buffered_input), .b(12'b001111011010), .eq(weq986));
    equaln #(12) e987(.a(buffered_input), .b(12'b001111011011), .eq(weq987));
    equaln #(12) e988(.a(buffered_input), .b(12'b001111011100), .eq(weq988));
    equaln #(12) e989(.a(buffered_input), .b(12'b001111011101), .eq(weq989));
    equaln #(12) e990(.a(buffered_input), .b(12'b001111011110), .eq(weq990));
    equaln #(12) e991(.a(buffered_input), .b(12'b001111011111), .eq(weq991));
    equaln #(12) e992(.a(buffered_input), .b(12'b001111100000), .eq(weq992));
    equaln #(12) e993(.a(buffered_input), .b(12'b001111100001), .eq(weq993));
    equaln #(12) e994(.a(buffered_input), .b(12'b001111100010), .eq(weq994));
    equaln #(12) e995(.a(buffered_input), .b(12'b001111100011), .eq(weq995));
    equaln #(12) e996(.a(buffered_input), .b(12'b001111100100), .eq(weq996));
    equaln #(12) e997(.a(buffered_input), .b(12'b001111100101), .eq(weq997));
    equaln #(12) e998(.a(buffered_input), .b(12'b001111100110), .eq(weq998));
    equaln #(12) e999(.a(buffered_input), .b(12'b001111100111), .eq(weq999));
    equaln #(12) e1000(.a(buffered_input), .b(12'b001111101000), .eq(weq1000));
    equaln #(12) e1001(.a(buffered_input), .b(12'b001111101001), .eq(weq1001));
    equaln #(12) e1002(.a(buffered_input), .b(12'b001111101010), .eq(weq1002));
    equaln #(12) e1003(.a(buffered_input), .b(12'b001111101011), .eq(weq1003));
    equaln #(12) e1004(.a(buffered_input), .b(12'b001111101100), .eq(weq1004));
    equaln #(12) e1005(.a(buffered_input), .b(12'b001111101101), .eq(weq1005));
    equaln #(12) e1006(.a(buffered_input), .b(12'b001111101110), .eq(weq1006));
    equaln #(12) e1007(.a(buffered_input), .b(12'b001111101111), .eq(weq1007));
    equaln #(12) e1008(.a(buffered_input), .b(12'b001111110000), .eq(weq1008));
    equaln #(12) e1009(.a(buffered_input), .b(12'b001111110001), .eq(weq1009));
    equaln #(12) e1010(.a(buffered_input), .b(12'b001111110010), .eq(weq1010));
    equaln #(12) e1011(.a(buffered_input), .b(12'b001111110011), .eq(weq1011));
    equaln #(12) e1012(.a(buffered_input), .b(12'b001111110100), .eq(weq1012));
    equaln #(12) e1013(.a(buffered_input), .b(12'b001111110101), .eq(weq1013));
    equaln #(12) e1014(.a(buffered_input), .b(12'b001111110110), .eq(weq1014));
    equaln #(12) e1015(.a(buffered_input), .b(12'b001111110111), .eq(weq1015));
    equaln #(12) e1016(.a(buffered_input), .b(12'b001111111000), .eq(weq1016));
    equaln #(12) e1017(.a(buffered_input), .b(12'b001111111001), .eq(weq1017));
    equaln #(12) e1018(.a(buffered_input), .b(12'b001111111010), .eq(weq1018));
    equaln #(12) e1019(.a(buffered_input), .b(12'b001111111011), .eq(weq1019));
    equaln #(12) e1020(.a(buffered_input), .b(12'b001111111100), .eq(weq1020));
    equaln #(12) e1021(.a(buffered_input), .b(12'b001111111101), .eq(weq1021));
    equaln #(12) e1022(.a(buffered_input), .b(12'b001111111110), .eq(weq1022));
    equaln #(12) e1023(.a(buffered_input), .b(12'b001111111111), .eq(weq1023));
    equaln #(12) e1024(.a(buffered_input), .b(12'b010000000000), .eq(weq1024));
    equaln #(12) e1025(.a(buffered_input), .b(12'b010000000001), .eq(weq1025));
    equaln #(12) e1026(.a(buffered_input), .b(12'b010000000010), .eq(weq1026));
    equaln #(12) e1027(.a(buffered_input), .b(12'b010000000011), .eq(weq1027));
    equaln #(12) e1028(.a(buffered_input), .b(12'b010000000100), .eq(weq1028));
    equaln #(12) e1029(.a(buffered_input), .b(12'b010000000101), .eq(weq1029));
    equaln #(12) e1030(.a(buffered_input), .b(12'b010000000110), .eq(weq1030));
    equaln #(12) e1031(.a(buffered_input), .b(12'b010000000111), .eq(weq1031));
    equaln #(12) e1032(.a(buffered_input), .b(12'b010000001000), .eq(weq1032));
    equaln #(12) e1033(.a(buffered_input), .b(12'b010000001001), .eq(weq1033));
    equaln #(12) e1034(.a(buffered_input), .b(12'b010000001010), .eq(weq1034));
    equaln #(12) e1035(.a(buffered_input), .b(12'b010000001011), .eq(weq1035));
    equaln #(12) e1036(.a(buffered_input), .b(12'b010000001100), .eq(weq1036));
    equaln #(12) e1037(.a(buffered_input), .b(12'b010000001101), .eq(weq1037));
    equaln #(12) e1038(.a(buffered_input), .b(12'b010000001110), .eq(weq1038));
    equaln #(12) e1039(.a(buffered_input), .b(12'b010000001111), .eq(weq1039));
    equaln #(12) e1040(.a(buffered_input), .b(12'b010000010000), .eq(weq1040));
    equaln #(12) e1041(.a(buffered_input), .b(12'b010000010001), .eq(weq1041));
    equaln #(12) e1042(.a(buffered_input), .b(12'b010000010010), .eq(weq1042));
    equaln #(12) e1043(.a(buffered_input), .b(12'b010000010011), .eq(weq1043));
    equaln #(12) e1044(.a(buffered_input), .b(12'b010000010100), .eq(weq1044));
    equaln #(12) e1045(.a(buffered_input), .b(12'b010000010101), .eq(weq1045));
    equaln #(12) e1046(.a(buffered_input), .b(12'b010000010110), .eq(weq1046));
    equaln #(12) e1047(.a(buffered_input), .b(12'b010000010111), .eq(weq1047));
    equaln #(12) e1048(.a(buffered_input), .b(12'b010000011000), .eq(weq1048));
    equaln #(12) e1049(.a(buffered_input), .b(12'b010000011001), .eq(weq1049));
    equaln #(12) e1050(.a(buffered_input), .b(12'b010000011010), .eq(weq1050));
    equaln #(12) e1051(.a(buffered_input), .b(12'b010000011011), .eq(weq1051));
    equaln #(12) e1052(.a(buffered_input), .b(12'b010000011100), .eq(weq1052));
    equaln #(12) e1053(.a(buffered_input), .b(12'b010000011101), .eq(weq1053));
    equaln #(12) e1054(.a(buffered_input), .b(12'b010000011110), .eq(weq1054));
    equaln #(12) e1055(.a(buffered_input), .b(12'b010000011111), .eq(weq1055));
    equaln #(12) e1056(.a(buffered_input), .b(12'b010000100000), .eq(weq1056));
    equaln #(12) e1057(.a(buffered_input), .b(12'b010000100001), .eq(weq1057));
    equaln #(12) e1058(.a(buffered_input), .b(12'b010000100010), .eq(weq1058));
    equaln #(12) e1059(.a(buffered_input), .b(12'b010000100011), .eq(weq1059));
    equaln #(12) e1060(.a(buffered_input), .b(12'b010000100100), .eq(weq1060));
    equaln #(12) e1061(.a(buffered_input), .b(12'b010000100101), .eq(weq1061));
    equaln #(12) e1062(.a(buffered_input), .b(12'b010000100110), .eq(weq1062));
    equaln #(12) e1063(.a(buffered_input), .b(12'b010000100111), .eq(weq1063));
    equaln #(12) e1064(.a(buffered_input), .b(12'b010000101000), .eq(weq1064));
    equaln #(12) e1065(.a(buffered_input), .b(12'b010000101001), .eq(weq1065));
    equaln #(12) e1066(.a(buffered_input), .b(12'b010000101010), .eq(weq1066));
    equaln #(12) e1067(.a(buffered_input), .b(12'b010000101011), .eq(weq1067));
    equaln #(12) e1068(.a(buffered_input), .b(12'b010000101100), .eq(weq1068));
    equaln #(12) e1069(.a(buffered_input), .b(12'b010000101101), .eq(weq1069));
    equaln #(12) e1070(.a(buffered_input), .b(12'b010000101110), .eq(weq1070));
    equaln #(12) e1071(.a(buffered_input), .b(12'b010000101111), .eq(weq1071));
    equaln #(12) e1072(.a(buffered_input), .b(12'b010000110000), .eq(weq1072));
    equaln #(12) e1073(.a(buffered_input), .b(12'b010000110001), .eq(weq1073));
    equaln #(12) e1074(.a(buffered_input), .b(12'b010000110010), .eq(weq1074));
    equaln #(12) e1075(.a(buffered_input), .b(12'b010000110011), .eq(weq1075));
    equaln #(12) e1076(.a(buffered_input), .b(12'b010000110100), .eq(weq1076));
    equaln #(12) e1077(.a(buffered_input), .b(12'b010000110101), .eq(weq1077));
    equaln #(12) e1078(.a(buffered_input), .b(12'b010000110110), .eq(weq1078));
    equaln #(12) e1079(.a(buffered_input), .b(12'b010000110111), .eq(weq1079));
    equaln #(12) e1080(.a(buffered_input), .b(12'b010000111000), .eq(weq1080));
    equaln #(12) e1081(.a(buffered_input), .b(12'b010000111001), .eq(weq1081));
    equaln #(12) e1082(.a(buffered_input), .b(12'b010000111010), .eq(weq1082));
    equaln #(12) e1083(.a(buffered_input), .b(12'b010000111011), .eq(weq1083));
    equaln #(12) e1084(.a(buffered_input), .b(12'b010000111100), .eq(weq1084));
    equaln #(12) e1085(.a(buffered_input), .b(12'b010000111101), .eq(weq1085));
    equaln #(12) e1086(.a(buffered_input), .b(12'b010000111110), .eq(weq1086));
    equaln #(12) e1087(.a(buffered_input), .b(12'b010000111111), .eq(weq1087));
    equaln #(12) e1088(.a(buffered_input), .b(12'b010001000000), .eq(weq1088));
    equaln #(12) e1089(.a(buffered_input), .b(12'b010001000001), .eq(weq1089));
    equaln #(12) e1090(.a(buffered_input), .b(12'b010001000010), .eq(weq1090));
    equaln #(12) e1091(.a(buffered_input), .b(12'b010001000011), .eq(weq1091));
    equaln #(12) e1092(.a(buffered_input), .b(12'b010001000100), .eq(weq1092));
    equaln #(12) e1093(.a(buffered_input), .b(12'b010001000101), .eq(weq1093));
    equaln #(12) e1094(.a(buffered_input), .b(12'b010001000110), .eq(weq1094));
    equaln #(12) e1095(.a(buffered_input), .b(12'b010001000111), .eq(weq1095));
    equaln #(12) e1096(.a(buffered_input), .b(12'b010001001000), .eq(weq1096));
    equaln #(12) e1097(.a(buffered_input), .b(12'b010001001001), .eq(weq1097));
    equaln #(12) e1098(.a(buffered_input), .b(12'b010001001010), .eq(weq1098));
    equaln #(12) e1099(.a(buffered_input), .b(12'b010001001011), .eq(weq1099));
    equaln #(12) e1100(.a(buffered_input), .b(12'b010001001100), .eq(weq1100));
    equaln #(12) e1101(.a(buffered_input), .b(12'b010001001101), .eq(weq1101));
    equaln #(12) e1102(.a(buffered_input), .b(12'b010001001110), .eq(weq1102));
    equaln #(12) e1103(.a(buffered_input), .b(12'b010001001111), .eq(weq1103));
    equaln #(12) e1104(.a(buffered_input), .b(12'b010001010000), .eq(weq1104));
    equaln #(12) e1105(.a(buffered_input), .b(12'b010001010001), .eq(weq1105));
    equaln #(12) e1106(.a(buffered_input), .b(12'b010001010010), .eq(weq1106));
    equaln #(12) e1107(.a(buffered_input), .b(12'b010001010011), .eq(weq1107));
    equaln #(12) e1108(.a(buffered_input), .b(12'b010001010100), .eq(weq1108));
    equaln #(12) e1109(.a(buffered_input), .b(12'b010001010101), .eq(weq1109));
    equaln #(12) e1110(.a(buffered_input), .b(12'b010001010110), .eq(weq1110));
    equaln #(12) e1111(.a(buffered_input), .b(12'b010001010111), .eq(weq1111));
    equaln #(12) e1112(.a(buffered_input), .b(12'b010001011000), .eq(weq1112));
    equaln #(12) e1113(.a(buffered_input), .b(12'b010001011001), .eq(weq1113));
    equaln #(12) e1114(.a(buffered_input), .b(12'b010001011010), .eq(weq1114));
    equaln #(12) e1115(.a(buffered_input), .b(12'b010001011011), .eq(weq1115));
    equaln #(12) e1116(.a(buffered_input), .b(12'b010001011100), .eq(weq1116));
    equaln #(12) e1117(.a(buffered_input), .b(12'b010001011101), .eq(weq1117));
    equaln #(12) e1118(.a(buffered_input), .b(12'b010001011110), .eq(weq1118));
    equaln #(12) e1119(.a(buffered_input), .b(12'b010001011111), .eq(weq1119));
    equaln #(12) e1120(.a(buffered_input), .b(12'b010001100000), .eq(weq1120));
    equaln #(12) e1121(.a(buffered_input), .b(12'b010001100001), .eq(weq1121));
    equaln #(12) e1122(.a(buffered_input), .b(12'b010001100010), .eq(weq1122));
    equaln #(12) e1123(.a(buffered_input), .b(12'b010001100011), .eq(weq1123));
    equaln #(12) e1124(.a(buffered_input), .b(12'b010001100100), .eq(weq1124));
    equaln #(12) e1125(.a(buffered_input), .b(12'b010001100101), .eq(weq1125));
    equaln #(12) e1126(.a(buffered_input), .b(12'b010001100110), .eq(weq1126));
    equaln #(12) e1127(.a(buffered_input), .b(12'b010001100111), .eq(weq1127));
    equaln #(12) e1128(.a(buffered_input), .b(12'b010001101000), .eq(weq1128));
    equaln #(12) e1129(.a(buffered_input), .b(12'b010001101001), .eq(weq1129));
    equaln #(12) e1130(.a(buffered_input), .b(12'b010001101010), .eq(weq1130));
    equaln #(12) e1131(.a(buffered_input), .b(12'b010001101011), .eq(weq1131));
    equaln #(12) e1132(.a(buffered_input), .b(12'b010001101100), .eq(weq1132));
    equaln #(12) e1133(.a(buffered_input), .b(12'b010001101101), .eq(weq1133));
    equaln #(12) e1134(.a(buffered_input), .b(12'b010001101110), .eq(weq1134));
    equaln #(12) e1135(.a(buffered_input), .b(12'b010001101111), .eq(weq1135));
    equaln #(12) e1136(.a(buffered_input), .b(12'b010001110000), .eq(weq1136));
    equaln #(12) e1137(.a(buffered_input), .b(12'b010001110001), .eq(weq1137));
    equaln #(12) e1138(.a(buffered_input), .b(12'b010001110010), .eq(weq1138));
    equaln #(12) e1139(.a(buffered_input), .b(12'b010001110011), .eq(weq1139));
    equaln #(12) e1140(.a(buffered_input), .b(12'b010001110100), .eq(weq1140));
    equaln #(12) e1141(.a(buffered_input), .b(12'b010001110101), .eq(weq1141));
    equaln #(12) e1142(.a(buffered_input), .b(12'b010001110110), .eq(weq1142));
    equaln #(12) e1143(.a(buffered_input), .b(12'b010001110111), .eq(weq1143));
    equaln #(12) e1144(.a(buffered_input), .b(12'b010001111000), .eq(weq1144));
    equaln #(12) e1145(.a(buffered_input), .b(12'b010001111001), .eq(weq1145));
    equaln #(12) e1146(.a(buffered_input), .b(12'b010001111010), .eq(weq1146));
    equaln #(12) e1147(.a(buffered_input), .b(12'b010001111011), .eq(weq1147));
    equaln #(12) e1148(.a(buffered_input), .b(12'b010001111100), .eq(weq1148));
    equaln #(12) e1149(.a(buffered_input), .b(12'b010001111101), .eq(weq1149));
    equaln #(12) e1150(.a(buffered_input), .b(12'b010001111110), .eq(weq1150));
    equaln #(12) e1151(.a(buffered_input), .b(12'b010001111111), .eq(weq1151));
    equaln #(12) e1152(.a(buffered_input), .b(12'b010010000000), .eq(weq1152));
    equaln #(12) e1153(.a(buffered_input), .b(12'b010010000001), .eq(weq1153));
    equaln #(12) e1154(.a(buffered_input), .b(12'b010010000010), .eq(weq1154));
    equaln #(12) e1155(.a(buffered_input), .b(12'b010010000011), .eq(weq1155));
    equaln #(12) e1156(.a(buffered_input), .b(12'b010010000100), .eq(weq1156));
    equaln #(12) e1157(.a(buffered_input), .b(12'b010010000101), .eq(weq1157));
    equaln #(12) e1158(.a(buffered_input), .b(12'b010010000110), .eq(weq1158));
    equaln #(12) e1159(.a(buffered_input), .b(12'b010010000111), .eq(weq1159));
    equaln #(12) e1160(.a(buffered_input), .b(12'b010010001000), .eq(weq1160));
    equaln #(12) e1161(.a(buffered_input), .b(12'b010010001001), .eq(weq1161));
    equaln #(12) e1162(.a(buffered_input), .b(12'b010010001010), .eq(weq1162));
    equaln #(12) e1163(.a(buffered_input), .b(12'b010010001011), .eq(weq1163));
    equaln #(12) e1164(.a(buffered_input), .b(12'b010010001100), .eq(weq1164));
    equaln #(12) e1165(.a(buffered_input), .b(12'b010010001101), .eq(weq1165));
    equaln #(12) e1166(.a(buffered_input), .b(12'b010010001110), .eq(weq1166));
    equaln #(12) e1167(.a(buffered_input), .b(12'b010010001111), .eq(weq1167));
    equaln #(12) e1168(.a(buffered_input), .b(12'b010010010000), .eq(weq1168));
    equaln #(12) e1169(.a(buffered_input), .b(12'b010010010001), .eq(weq1169));
    equaln #(12) e1170(.a(buffered_input), .b(12'b010010010010), .eq(weq1170));
    equaln #(12) e1171(.a(buffered_input), .b(12'b010010010011), .eq(weq1171));
    equaln #(12) e1172(.a(buffered_input), .b(12'b010010010100), .eq(weq1172));
    equaln #(12) e1173(.a(buffered_input), .b(12'b010010010101), .eq(weq1173));
    equaln #(12) e1174(.a(buffered_input), .b(12'b010010010110), .eq(weq1174));
    equaln #(12) e1175(.a(buffered_input), .b(12'b010010010111), .eq(weq1175));
    equaln #(12) e1176(.a(buffered_input), .b(12'b010010011000), .eq(weq1176));
    equaln #(12) e1177(.a(buffered_input), .b(12'b010010011001), .eq(weq1177));
    equaln #(12) e1178(.a(buffered_input), .b(12'b010010011010), .eq(weq1178));
    equaln #(12) e1179(.a(buffered_input), .b(12'b010010011011), .eq(weq1179));
    equaln #(12) e1180(.a(buffered_input), .b(12'b010010011100), .eq(weq1180));
    equaln #(12) e1181(.a(buffered_input), .b(12'b010010011101), .eq(weq1181));
    equaln #(12) e1182(.a(buffered_input), .b(12'b010010011110), .eq(weq1182));
    equaln #(12) e1183(.a(buffered_input), .b(12'b010010011111), .eq(weq1183));
    equaln #(12) e1184(.a(buffered_input), .b(12'b010010100000), .eq(weq1184));
    equaln #(12) e1185(.a(buffered_input), .b(12'b010010100001), .eq(weq1185));
    equaln #(12) e1186(.a(buffered_input), .b(12'b010010100010), .eq(weq1186));
    equaln #(12) e1187(.a(buffered_input), .b(12'b010010100011), .eq(weq1187));
    equaln #(12) e1188(.a(buffered_input), .b(12'b010010100100), .eq(weq1188));
    equaln #(12) e1189(.a(buffered_input), .b(12'b010010100101), .eq(weq1189));
    equaln #(12) e1190(.a(buffered_input), .b(12'b010010100110), .eq(weq1190));
    equaln #(12) e1191(.a(buffered_input), .b(12'b010010100111), .eq(weq1191));
    equaln #(12) e1192(.a(buffered_input), .b(12'b010010101000), .eq(weq1192));
    equaln #(12) e1193(.a(buffered_input), .b(12'b010010101001), .eq(weq1193));
    equaln #(12) e1194(.a(buffered_input), .b(12'b010010101010), .eq(weq1194));
    equaln #(12) e1195(.a(buffered_input), .b(12'b010010101011), .eq(weq1195));
    equaln #(12) e1196(.a(buffered_input), .b(12'b010010101100), .eq(weq1196));
    equaln #(12) e1197(.a(buffered_input), .b(12'b010010101101), .eq(weq1197));
    equaln #(12) e1198(.a(buffered_input), .b(12'b010010101110), .eq(weq1198));
    equaln #(12) e1199(.a(buffered_input), .b(12'b010010101111), .eq(weq1199));
    equaln #(12) e1200(.a(buffered_input), .b(12'b010010110000), .eq(weq1200));
    equaln #(12) e1201(.a(buffered_input), .b(12'b010010110001), .eq(weq1201));
    equaln #(12) e1202(.a(buffered_input), .b(12'b010010110010), .eq(weq1202));
    equaln #(12) e1203(.a(buffered_input), .b(12'b010010110011), .eq(weq1203));
    equaln #(12) e1204(.a(buffered_input), .b(12'b010010110100), .eq(weq1204));
    equaln #(12) e1205(.a(buffered_input), .b(12'b010010110101), .eq(weq1205));
    equaln #(12) e1206(.a(buffered_input), .b(12'b010010110110), .eq(weq1206));
    equaln #(12) e1207(.a(buffered_input), .b(12'b010010110111), .eq(weq1207));
    equaln #(12) e1208(.a(buffered_input), .b(12'b010010111000), .eq(weq1208));
    equaln #(12) e1209(.a(buffered_input), .b(12'b010010111001), .eq(weq1209));
    equaln #(12) e1210(.a(buffered_input), .b(12'b010010111010), .eq(weq1210));
    equaln #(12) e1211(.a(buffered_input), .b(12'b010010111011), .eq(weq1211));
    equaln #(12) e1212(.a(buffered_input), .b(12'b010010111100), .eq(weq1212));
    equaln #(12) e1213(.a(buffered_input), .b(12'b010010111101), .eq(weq1213));
    equaln #(12) e1214(.a(buffered_input), .b(12'b010010111110), .eq(weq1214));
    equaln #(12) e1215(.a(buffered_input), .b(12'b010010111111), .eq(weq1215));
    equaln #(12) e1216(.a(buffered_input), .b(12'b010011000000), .eq(weq1216));
    equaln #(12) e1217(.a(buffered_input), .b(12'b010011000001), .eq(weq1217));
    equaln #(12) e1218(.a(buffered_input), .b(12'b010011000010), .eq(weq1218));
    equaln #(12) e1219(.a(buffered_input), .b(12'b010011000011), .eq(weq1219));
    equaln #(12) e1220(.a(buffered_input), .b(12'b010011000100), .eq(weq1220));
    equaln #(12) e1221(.a(buffered_input), .b(12'b010011000101), .eq(weq1221));
    equaln #(12) e1222(.a(buffered_input), .b(12'b010011000110), .eq(weq1222));
    equaln #(12) e1223(.a(buffered_input), .b(12'b010011000111), .eq(weq1223));
    equaln #(12) e1224(.a(buffered_input), .b(12'b010011001000), .eq(weq1224));
    equaln #(12) e1225(.a(buffered_input), .b(12'b010011001001), .eq(weq1225));
    equaln #(12) e1226(.a(buffered_input), .b(12'b010011001010), .eq(weq1226));
    equaln #(12) e1227(.a(buffered_input), .b(12'b010011001011), .eq(weq1227));
    equaln #(12) e1228(.a(buffered_input), .b(12'b010011001100), .eq(weq1228));
    equaln #(12) e1229(.a(buffered_input), .b(12'b010011001101), .eq(weq1229));
    equaln #(12) e1230(.a(buffered_input), .b(12'b010011001110), .eq(weq1230));
    equaln #(12) e1231(.a(buffered_input), .b(12'b010011001111), .eq(weq1231));
    equaln #(12) e1232(.a(buffered_input), .b(12'b010011010000), .eq(weq1232));
    equaln #(12) e1233(.a(buffered_input), .b(12'b010011010001), .eq(weq1233));
    equaln #(12) e1234(.a(buffered_input), .b(12'b010011010010), .eq(weq1234));
    equaln #(12) e1235(.a(buffered_input), .b(12'b010011010011), .eq(weq1235));
    equaln #(12) e1236(.a(buffered_input), .b(12'b010011010100), .eq(weq1236));
    equaln #(12) e1237(.a(buffered_input), .b(12'b010011010101), .eq(weq1237));
    equaln #(12) e1238(.a(buffered_input), .b(12'b010011010110), .eq(weq1238));
    equaln #(12) e1239(.a(buffered_input), .b(12'b010011010111), .eq(weq1239));
    equaln #(12) e1240(.a(buffered_input), .b(12'b010011011000), .eq(weq1240));
    equaln #(12) e1241(.a(buffered_input), .b(12'b010011011001), .eq(weq1241));
    equaln #(12) e1242(.a(buffered_input), .b(12'b010011011010), .eq(weq1242));
    equaln #(12) e1243(.a(buffered_input), .b(12'b010011011011), .eq(weq1243));
    equaln #(12) e1244(.a(buffered_input), .b(12'b010011011100), .eq(weq1244));
    equaln #(12) e1245(.a(buffered_input), .b(12'b010011011101), .eq(weq1245));
    equaln #(12) e1246(.a(buffered_input), .b(12'b010011011110), .eq(weq1246));
    equaln #(12) e1247(.a(buffered_input), .b(12'b010011011111), .eq(weq1247));
    equaln #(12) e1248(.a(buffered_input), .b(12'b010011100000), .eq(weq1248));
    equaln #(12) e1249(.a(buffered_input), .b(12'b010011100001), .eq(weq1249));
    equaln #(12) e1250(.a(buffered_input), .b(12'b010011100010), .eq(weq1250));
    equaln #(12) e1251(.a(buffered_input), .b(12'b010011100011), .eq(weq1251));
    equaln #(12) e1252(.a(buffered_input), .b(12'b010011100100), .eq(weq1252));
    equaln #(12) e1253(.a(buffered_input), .b(12'b010011100101), .eq(weq1253));
    equaln #(12) e1254(.a(buffered_input), .b(12'b010011100110), .eq(weq1254));
    equaln #(12) e1255(.a(buffered_input), .b(12'b010011100111), .eq(weq1255));
    equaln #(12) e1256(.a(buffered_input), .b(12'b010011101000), .eq(weq1256));
    equaln #(12) e1257(.a(buffered_input), .b(12'b010011101001), .eq(weq1257));
    equaln #(12) e1258(.a(buffered_input), .b(12'b010011101010), .eq(weq1258));
    equaln #(12) e1259(.a(buffered_input), .b(12'b010011101011), .eq(weq1259));
    equaln #(12) e1260(.a(buffered_input), .b(12'b010011101100), .eq(weq1260));
    equaln #(12) e1261(.a(buffered_input), .b(12'b010011101101), .eq(weq1261));
    equaln #(12) e1262(.a(buffered_input), .b(12'b010011101110), .eq(weq1262));
    equaln #(12) e1263(.a(buffered_input), .b(12'b010011101111), .eq(weq1263));
    equaln #(12) e1264(.a(buffered_input), .b(12'b010011110000), .eq(weq1264));
    equaln #(12) e1265(.a(buffered_input), .b(12'b010011110001), .eq(weq1265));
    equaln #(12) e1266(.a(buffered_input), .b(12'b010011110010), .eq(weq1266));
    equaln #(12) e1267(.a(buffered_input), .b(12'b010011110011), .eq(weq1267));
    equaln #(12) e1268(.a(buffered_input), .b(12'b010011110100), .eq(weq1268));
    equaln #(12) e1269(.a(buffered_input), .b(12'b010011110101), .eq(weq1269));
    equaln #(12) e1270(.a(buffered_input), .b(12'b010011110110), .eq(weq1270));
    equaln #(12) e1271(.a(buffered_input), .b(12'b010011110111), .eq(weq1271));
    equaln #(12) e1272(.a(buffered_input), .b(12'b010011111000), .eq(weq1272));
    equaln #(12) e1273(.a(buffered_input), .b(12'b010011111001), .eq(weq1273));
    equaln #(12) e1274(.a(buffered_input), .b(12'b010011111010), .eq(weq1274));
    equaln #(12) e1275(.a(buffered_input), .b(12'b010011111011), .eq(weq1275));
    equaln #(12) e1276(.a(buffered_input), .b(12'b010011111100), .eq(weq1276));
    equaln #(12) e1277(.a(buffered_input), .b(12'b010011111101), .eq(weq1277));
    equaln #(12) e1278(.a(buffered_input), .b(12'b010011111110), .eq(weq1278));
    equaln #(12) e1279(.a(buffered_input), .b(12'b010011111111), .eq(weq1279));
    equaln #(12) e1280(.a(buffered_input), .b(12'b010100000000), .eq(weq1280));
    equaln #(12) e1281(.a(buffered_input), .b(12'b010100000001), .eq(weq1281));
    equaln #(12) e1282(.a(buffered_input), .b(12'b010100000010), .eq(weq1282));
    equaln #(12) e1283(.a(buffered_input), .b(12'b010100000011), .eq(weq1283));
    equaln #(12) e1284(.a(buffered_input), .b(12'b010100000100), .eq(weq1284));
    equaln #(12) e1285(.a(buffered_input), .b(12'b010100000101), .eq(weq1285));
    equaln #(12) e1286(.a(buffered_input), .b(12'b010100000110), .eq(weq1286));
    equaln #(12) e1287(.a(buffered_input), .b(12'b010100000111), .eq(weq1287));
    equaln #(12) e1288(.a(buffered_input), .b(12'b010100001000), .eq(weq1288));
    equaln #(12) e1289(.a(buffered_input), .b(12'b010100001001), .eq(weq1289));
    equaln #(12) e1290(.a(buffered_input), .b(12'b010100001010), .eq(weq1290));
    equaln #(12) e1291(.a(buffered_input), .b(12'b010100001011), .eq(weq1291));
    equaln #(12) e1292(.a(buffered_input), .b(12'b010100001100), .eq(weq1292));
    equaln #(12) e1293(.a(buffered_input), .b(12'b010100001101), .eq(weq1293));
    equaln #(12) e1294(.a(buffered_input), .b(12'b010100001110), .eq(weq1294));
    equaln #(12) e1295(.a(buffered_input), .b(12'b010100001111), .eq(weq1295));
    equaln #(12) e1296(.a(buffered_input), .b(12'b010100010000), .eq(weq1296));
    equaln #(12) e1297(.a(buffered_input), .b(12'b010100010001), .eq(weq1297));
    equaln #(12) e1298(.a(buffered_input), .b(12'b010100010010), .eq(weq1298));
    equaln #(12) e1299(.a(buffered_input), .b(12'b010100010011), .eq(weq1299));
    equaln #(12) e1300(.a(buffered_input), .b(12'b010100010100), .eq(weq1300));
    equaln #(12) e1301(.a(buffered_input), .b(12'b010100010101), .eq(weq1301));
    equaln #(12) e1302(.a(buffered_input), .b(12'b010100010110), .eq(weq1302));
    equaln #(12) e1303(.a(buffered_input), .b(12'b010100010111), .eq(weq1303));
    equaln #(12) e1304(.a(buffered_input), .b(12'b010100011000), .eq(weq1304));
    equaln #(12) e1305(.a(buffered_input), .b(12'b010100011001), .eq(weq1305));
    equaln #(12) e1306(.a(buffered_input), .b(12'b010100011010), .eq(weq1306));
    equaln #(12) e1307(.a(buffered_input), .b(12'b010100011011), .eq(weq1307));
    equaln #(12) e1308(.a(buffered_input), .b(12'b010100011100), .eq(weq1308));
    equaln #(12) e1309(.a(buffered_input), .b(12'b010100011101), .eq(weq1309));
    equaln #(12) e1310(.a(buffered_input), .b(12'b010100011110), .eq(weq1310));
    equaln #(12) e1311(.a(buffered_input), .b(12'b010100011111), .eq(weq1311));
    equaln #(12) e1312(.a(buffered_input), .b(12'b010100100000), .eq(weq1312));
    equaln #(12) e1313(.a(buffered_input), .b(12'b010100100001), .eq(weq1313));
    equaln #(12) e1314(.a(buffered_input), .b(12'b010100100010), .eq(weq1314));
    equaln #(12) e1315(.a(buffered_input), .b(12'b010100100011), .eq(weq1315));
    equaln #(12) e1316(.a(buffered_input), .b(12'b010100100100), .eq(weq1316));
    equaln #(12) e1317(.a(buffered_input), .b(12'b010100100101), .eq(weq1317));
    equaln #(12) e1318(.a(buffered_input), .b(12'b010100100110), .eq(weq1318));
    equaln #(12) e1319(.a(buffered_input), .b(12'b010100100111), .eq(weq1319));
    equaln #(12) e1320(.a(buffered_input), .b(12'b010100101000), .eq(weq1320));
    equaln #(12) e1321(.a(buffered_input), .b(12'b010100101001), .eq(weq1321));
    equaln #(12) e1322(.a(buffered_input), .b(12'b010100101010), .eq(weq1322));
    equaln #(12) e1323(.a(buffered_input), .b(12'b010100101011), .eq(weq1323));
    equaln #(12) e1324(.a(buffered_input), .b(12'b010100101100), .eq(weq1324));
    equaln #(12) e1325(.a(buffered_input), .b(12'b010100101101), .eq(weq1325));
    equaln #(12) e1326(.a(buffered_input), .b(12'b010100101110), .eq(weq1326));
    equaln #(12) e1327(.a(buffered_input), .b(12'b010100101111), .eq(weq1327));
    equaln #(12) e1328(.a(buffered_input), .b(12'b010100110000), .eq(weq1328));
    equaln #(12) e1329(.a(buffered_input), .b(12'b010100110001), .eq(weq1329));
    equaln #(12) e1330(.a(buffered_input), .b(12'b010100110010), .eq(weq1330));
    equaln #(12) e1331(.a(buffered_input), .b(12'b010100110011), .eq(weq1331));
    equaln #(12) e1332(.a(buffered_input), .b(12'b010100110100), .eq(weq1332));
    equaln #(12) e1333(.a(buffered_input), .b(12'b010100110101), .eq(weq1333));
    equaln #(12) e1334(.a(buffered_input), .b(12'b010100110110), .eq(weq1334));
    equaln #(12) e1335(.a(buffered_input), .b(12'b010100110111), .eq(weq1335));
    equaln #(12) e1336(.a(buffered_input), .b(12'b010100111000), .eq(weq1336));
    equaln #(12) e1337(.a(buffered_input), .b(12'b010100111001), .eq(weq1337));
    equaln #(12) e1338(.a(buffered_input), .b(12'b010100111010), .eq(weq1338));
    equaln #(12) e1339(.a(buffered_input), .b(12'b010100111011), .eq(weq1339));
    equaln #(12) e1340(.a(buffered_input), .b(12'b010100111100), .eq(weq1340));
    equaln #(12) e1341(.a(buffered_input), .b(12'b010100111101), .eq(weq1341));
    equaln #(12) e1342(.a(buffered_input), .b(12'b010100111110), .eq(weq1342));
    equaln #(12) e1343(.a(buffered_input), .b(12'b010100111111), .eq(weq1343));
    equaln #(12) e1344(.a(buffered_input), .b(12'b010101000000), .eq(weq1344));
    equaln #(12) e1345(.a(buffered_input), .b(12'b010101000001), .eq(weq1345));
    equaln #(12) e1346(.a(buffered_input), .b(12'b010101000010), .eq(weq1346));
    equaln #(12) e1347(.a(buffered_input), .b(12'b010101000011), .eq(weq1347));
    equaln #(12) e1348(.a(buffered_input), .b(12'b010101000100), .eq(weq1348));
    equaln #(12) e1349(.a(buffered_input), .b(12'b010101000101), .eq(weq1349));
    equaln #(12) e1350(.a(buffered_input), .b(12'b010101000110), .eq(weq1350));
    equaln #(12) e1351(.a(buffered_input), .b(12'b010101000111), .eq(weq1351));
    equaln #(12) e1352(.a(buffered_input), .b(12'b010101001000), .eq(weq1352));
    equaln #(12) e1353(.a(buffered_input), .b(12'b010101001001), .eq(weq1353));
    equaln #(12) e1354(.a(buffered_input), .b(12'b010101001010), .eq(weq1354));
    equaln #(12) e1355(.a(buffered_input), .b(12'b010101001011), .eq(weq1355));
    equaln #(12) e1356(.a(buffered_input), .b(12'b010101001100), .eq(weq1356));
    equaln #(12) e1357(.a(buffered_input), .b(12'b010101001101), .eq(weq1357));
    equaln #(12) e1358(.a(buffered_input), .b(12'b010101001110), .eq(weq1358));
    equaln #(12) e1359(.a(buffered_input), .b(12'b010101001111), .eq(weq1359));
    equaln #(12) e1360(.a(buffered_input), .b(12'b010101010000), .eq(weq1360));
    equaln #(12) e1361(.a(buffered_input), .b(12'b010101010001), .eq(weq1361));
    equaln #(12) e1362(.a(buffered_input), .b(12'b010101010010), .eq(weq1362));
    equaln #(12) e1363(.a(buffered_input), .b(12'b010101010011), .eq(weq1363));
    equaln #(12) e1364(.a(buffered_input), .b(12'b010101010100), .eq(weq1364));
    equaln #(12) e1365(.a(buffered_input), .b(12'b010101010101), .eq(weq1365));
    equaln #(12) e1366(.a(buffered_input), .b(12'b010101010110), .eq(weq1366));
    equaln #(12) e1367(.a(buffered_input), .b(12'b010101010111), .eq(weq1367));
    equaln #(12) e1368(.a(buffered_input), .b(12'b010101011000), .eq(weq1368));
    equaln #(12) e1369(.a(buffered_input), .b(12'b010101011001), .eq(weq1369));
    equaln #(12) e1370(.a(buffered_input), .b(12'b010101011010), .eq(weq1370));
    equaln #(12) e1371(.a(buffered_input), .b(12'b010101011011), .eq(weq1371));
    equaln #(12) e1372(.a(buffered_input), .b(12'b010101011100), .eq(weq1372));
    equaln #(12) e1373(.a(buffered_input), .b(12'b010101011101), .eq(weq1373));
    equaln #(12) e1374(.a(buffered_input), .b(12'b010101011110), .eq(weq1374));
    equaln #(12) e1375(.a(buffered_input), .b(12'b010101011111), .eq(weq1375));
    equaln #(12) e1376(.a(buffered_input), .b(12'b010101100000), .eq(weq1376));
    equaln #(12) e1377(.a(buffered_input), .b(12'b010101100001), .eq(weq1377));
    equaln #(12) e1378(.a(buffered_input), .b(12'b010101100010), .eq(weq1378));
    equaln #(12) e1379(.a(buffered_input), .b(12'b010101100011), .eq(weq1379));
    equaln #(12) e1380(.a(buffered_input), .b(12'b010101100100), .eq(weq1380));
    equaln #(12) e1381(.a(buffered_input), .b(12'b010101100101), .eq(weq1381));
    equaln #(12) e1382(.a(buffered_input), .b(12'b010101100110), .eq(weq1382));
    equaln #(12) e1383(.a(buffered_input), .b(12'b010101100111), .eq(weq1383));
    equaln #(12) e1384(.a(buffered_input), .b(12'b010101101000), .eq(weq1384));
    equaln #(12) e1385(.a(buffered_input), .b(12'b010101101001), .eq(weq1385));
    equaln #(12) e1386(.a(buffered_input), .b(12'b010101101010), .eq(weq1386));
    equaln #(12) e1387(.a(buffered_input), .b(12'b010101101011), .eq(weq1387));
    equaln #(12) e1388(.a(buffered_input), .b(12'b010101101100), .eq(weq1388));
    equaln #(12) e1389(.a(buffered_input), .b(12'b010101101101), .eq(weq1389));
    equaln #(12) e1390(.a(buffered_input), .b(12'b010101101110), .eq(weq1390));
    equaln #(12) e1391(.a(buffered_input), .b(12'b010101101111), .eq(weq1391));
    equaln #(12) e1392(.a(buffered_input), .b(12'b010101110000), .eq(weq1392));
    equaln #(12) e1393(.a(buffered_input), .b(12'b010101110001), .eq(weq1393));
    equaln #(12) e1394(.a(buffered_input), .b(12'b010101110010), .eq(weq1394));
    equaln #(12) e1395(.a(buffered_input), .b(12'b010101110011), .eq(weq1395));
    equaln #(12) e1396(.a(buffered_input), .b(12'b010101110100), .eq(weq1396));
    equaln #(12) e1397(.a(buffered_input), .b(12'b010101110101), .eq(weq1397));
    equaln #(12) e1398(.a(buffered_input), .b(12'b010101110110), .eq(weq1398));
    equaln #(12) e1399(.a(buffered_input), .b(12'b010101110111), .eq(weq1399));
    equaln #(12) e1400(.a(buffered_input), .b(12'b010101111000), .eq(weq1400));
    equaln #(12) e1401(.a(buffered_input), .b(12'b010101111001), .eq(weq1401));
    equaln #(12) e1402(.a(buffered_input), .b(12'b010101111010), .eq(weq1402));
    equaln #(12) e1403(.a(buffered_input), .b(12'b010101111011), .eq(weq1403));
    equaln #(12) e1404(.a(buffered_input), .b(12'b010101111100), .eq(weq1404));
    equaln #(12) e1405(.a(buffered_input), .b(12'b010101111101), .eq(weq1405));
    equaln #(12) e1406(.a(buffered_input), .b(12'b010101111110), .eq(weq1406));
    equaln #(12) e1407(.a(buffered_input), .b(12'b010101111111), .eq(weq1407));
    equaln #(12) e1408(.a(buffered_input), .b(12'b010110000000), .eq(weq1408));
    equaln #(12) e1409(.a(buffered_input), .b(12'b010110000001), .eq(weq1409));
    equaln #(12) e1410(.a(buffered_input), .b(12'b010110000010), .eq(weq1410));
    equaln #(12) e1411(.a(buffered_input), .b(12'b010110000011), .eq(weq1411));
    equaln #(12) e1412(.a(buffered_input), .b(12'b010110000100), .eq(weq1412));
    equaln #(12) e1413(.a(buffered_input), .b(12'b010110000101), .eq(weq1413));
    equaln #(12) e1414(.a(buffered_input), .b(12'b010110000110), .eq(weq1414));
    equaln #(12) e1415(.a(buffered_input), .b(12'b010110000111), .eq(weq1415));
    equaln #(12) e1416(.a(buffered_input), .b(12'b010110001000), .eq(weq1416));
    equaln #(12) e1417(.a(buffered_input), .b(12'b010110001001), .eq(weq1417));
    equaln #(12) e1418(.a(buffered_input), .b(12'b010110001010), .eq(weq1418));
    equaln #(12) e1419(.a(buffered_input), .b(12'b010110001011), .eq(weq1419));
    equaln #(12) e1420(.a(buffered_input), .b(12'b010110001100), .eq(weq1420));
    equaln #(12) e1421(.a(buffered_input), .b(12'b010110001101), .eq(weq1421));
    equaln #(12) e1422(.a(buffered_input), .b(12'b010110001110), .eq(weq1422));
    equaln #(12) e1423(.a(buffered_input), .b(12'b010110001111), .eq(weq1423));
    equaln #(12) e1424(.a(buffered_input), .b(12'b010110010000), .eq(weq1424));
    equaln #(12) e1425(.a(buffered_input), .b(12'b010110010001), .eq(weq1425));
    equaln #(12) e1426(.a(buffered_input), .b(12'b010110010010), .eq(weq1426));
    equaln #(12) e1427(.a(buffered_input), .b(12'b010110010011), .eq(weq1427));
    equaln #(12) e1428(.a(buffered_input), .b(12'b010110010100), .eq(weq1428));
    equaln #(12) e1429(.a(buffered_input), .b(12'b010110010101), .eq(weq1429));
    equaln #(12) e1430(.a(buffered_input), .b(12'b010110010110), .eq(weq1430));
    equaln #(12) e1431(.a(buffered_input), .b(12'b010110010111), .eq(weq1431));
    equaln #(12) e1432(.a(buffered_input), .b(12'b010110011000), .eq(weq1432));
    equaln #(12) e1433(.a(buffered_input), .b(12'b010110011001), .eq(weq1433));
    equaln #(12) e1434(.a(buffered_input), .b(12'b010110011010), .eq(weq1434));
    equaln #(12) e1435(.a(buffered_input), .b(12'b010110011011), .eq(weq1435));
    equaln #(12) e1436(.a(buffered_input), .b(12'b010110011100), .eq(weq1436));
    equaln #(12) e1437(.a(buffered_input), .b(12'b010110011101), .eq(weq1437));
    equaln #(12) e1438(.a(buffered_input), .b(12'b010110011110), .eq(weq1438));
    equaln #(12) e1439(.a(buffered_input), .b(12'b010110011111), .eq(weq1439));
    equaln #(12) e1440(.a(buffered_input), .b(12'b010110100000), .eq(weq1440));
    equaln #(12) e1441(.a(buffered_input), .b(12'b010110100001), .eq(weq1441));
    equaln #(12) e1442(.a(buffered_input), .b(12'b010110100010), .eq(weq1442));
    equaln #(12) e1443(.a(buffered_input), .b(12'b010110100011), .eq(weq1443));
    equaln #(12) e1444(.a(buffered_input), .b(12'b010110100100), .eq(weq1444));
    equaln #(12) e1445(.a(buffered_input), .b(12'b010110100101), .eq(weq1445));
    equaln #(12) e1446(.a(buffered_input), .b(12'b010110100110), .eq(weq1446));
    equaln #(12) e1447(.a(buffered_input), .b(12'b010110100111), .eq(weq1447));
    equaln #(12) e1448(.a(buffered_input), .b(12'b010110101000), .eq(weq1448));
    equaln #(12) e1449(.a(buffered_input), .b(12'b010110101001), .eq(weq1449));
    equaln #(12) e1450(.a(buffered_input), .b(12'b010110101010), .eq(weq1450));
    equaln #(12) e1451(.a(buffered_input), .b(12'b010110101011), .eq(weq1451));
    equaln #(12) e1452(.a(buffered_input), .b(12'b010110101100), .eq(weq1452));
    equaln #(12) e1453(.a(buffered_input), .b(12'b010110101101), .eq(weq1453));
    equaln #(12) e1454(.a(buffered_input), .b(12'b010110101110), .eq(weq1454));
    equaln #(12) e1455(.a(buffered_input), .b(12'b010110101111), .eq(weq1455));
    equaln #(12) e1456(.a(buffered_input), .b(12'b010110110000), .eq(weq1456));
    equaln #(12) e1457(.a(buffered_input), .b(12'b010110110001), .eq(weq1457));
    equaln #(12) e1458(.a(buffered_input), .b(12'b010110110010), .eq(weq1458));
    equaln #(12) e1459(.a(buffered_input), .b(12'b010110110011), .eq(weq1459));
    equaln #(12) e1460(.a(buffered_input), .b(12'b010110110100), .eq(weq1460));
    equaln #(12) e1461(.a(buffered_input), .b(12'b010110110101), .eq(weq1461));
    equaln #(12) e1462(.a(buffered_input), .b(12'b010110110110), .eq(weq1462));
    equaln #(12) e1463(.a(buffered_input), .b(12'b010110110111), .eq(weq1463));
    equaln #(12) e1464(.a(buffered_input), .b(12'b010110111000), .eq(weq1464));
    equaln #(12) e1465(.a(buffered_input), .b(12'b010110111001), .eq(weq1465));
    equaln #(12) e1466(.a(buffered_input), .b(12'b010110111010), .eq(weq1466));
    equaln #(12) e1467(.a(buffered_input), .b(12'b010110111011), .eq(weq1467));
    equaln #(12) e1468(.a(buffered_input), .b(12'b010110111100), .eq(weq1468));
    equaln #(12) e1469(.a(buffered_input), .b(12'b010110111101), .eq(weq1469));
    equaln #(12) e1470(.a(buffered_input), .b(12'b010110111110), .eq(weq1470));
    equaln #(12) e1471(.a(buffered_input), .b(12'b010110111111), .eq(weq1471));
    equaln #(12) e1472(.a(buffered_input), .b(12'b010111000000), .eq(weq1472));
    equaln #(12) e1473(.a(buffered_input), .b(12'b010111000001), .eq(weq1473));
    equaln #(12) e1474(.a(buffered_input), .b(12'b010111000010), .eq(weq1474));
    equaln #(12) e1475(.a(buffered_input), .b(12'b010111000011), .eq(weq1475));
    equaln #(12) e1476(.a(buffered_input), .b(12'b010111000100), .eq(weq1476));
    equaln #(12) e1477(.a(buffered_input), .b(12'b010111000101), .eq(weq1477));
    equaln #(12) e1478(.a(buffered_input), .b(12'b010111000110), .eq(weq1478));
    equaln #(12) e1479(.a(buffered_input), .b(12'b010111000111), .eq(weq1479));
    equaln #(12) e1480(.a(buffered_input), .b(12'b010111001000), .eq(weq1480));
    equaln #(12) e1481(.a(buffered_input), .b(12'b010111001001), .eq(weq1481));
    equaln #(12) e1482(.a(buffered_input), .b(12'b010111001010), .eq(weq1482));
    equaln #(12) e1483(.a(buffered_input), .b(12'b010111001011), .eq(weq1483));
    equaln #(12) e1484(.a(buffered_input), .b(12'b010111001100), .eq(weq1484));
    equaln #(12) e1485(.a(buffered_input), .b(12'b010111001101), .eq(weq1485));
    equaln #(12) e1486(.a(buffered_input), .b(12'b010111001110), .eq(weq1486));
    equaln #(12) e1487(.a(buffered_input), .b(12'b010111001111), .eq(weq1487));
    equaln #(12) e1488(.a(buffered_input), .b(12'b010111010000), .eq(weq1488));
    equaln #(12) e1489(.a(buffered_input), .b(12'b010111010001), .eq(weq1489));
    equaln #(12) e1490(.a(buffered_input), .b(12'b010111010010), .eq(weq1490));
    equaln #(12) e1491(.a(buffered_input), .b(12'b010111010011), .eq(weq1491));
    equaln #(12) e1492(.a(buffered_input), .b(12'b010111010100), .eq(weq1492));
    equaln #(12) e1493(.a(buffered_input), .b(12'b010111010101), .eq(weq1493));
    equaln #(12) e1494(.a(buffered_input), .b(12'b010111010110), .eq(weq1494));
    equaln #(12) e1495(.a(buffered_input), .b(12'b010111010111), .eq(weq1495));
    equaln #(12) e1496(.a(buffered_input), .b(12'b010111011000), .eq(weq1496));
    equaln #(12) e1497(.a(buffered_input), .b(12'b010111011001), .eq(weq1497));
    equaln #(12) e1498(.a(buffered_input), .b(12'b010111011010), .eq(weq1498));
    equaln #(12) e1499(.a(buffered_input), .b(12'b010111011011), .eq(weq1499));
    equaln #(12) e1500(.a(buffered_input), .b(12'b010111011100), .eq(weq1500));
    equaln #(12) e1501(.a(buffered_input), .b(12'b010111011101), .eq(weq1501));
    equaln #(12) e1502(.a(buffered_input), .b(12'b010111011110), .eq(weq1502));
    equaln #(12) e1503(.a(buffered_input), .b(12'b010111011111), .eq(weq1503));
    equaln #(12) e1504(.a(buffered_input), .b(12'b010111100000), .eq(weq1504));
    equaln #(12) e1505(.a(buffered_input), .b(12'b010111100001), .eq(weq1505));
    equaln #(12) e1506(.a(buffered_input), .b(12'b010111100010), .eq(weq1506));
    equaln #(12) e1507(.a(buffered_input), .b(12'b010111100011), .eq(weq1507));
    equaln #(12) e1508(.a(buffered_input), .b(12'b010111100100), .eq(weq1508));
    equaln #(12) e1509(.a(buffered_input), .b(12'b010111100101), .eq(weq1509));
    equaln #(12) e1510(.a(buffered_input), .b(12'b010111100110), .eq(weq1510));
    equaln #(12) e1511(.a(buffered_input), .b(12'b010111100111), .eq(weq1511));
    equaln #(12) e1512(.a(buffered_input), .b(12'b010111101000), .eq(weq1512));
    equaln #(12) e1513(.a(buffered_input), .b(12'b010111101001), .eq(weq1513));
    equaln #(12) e1514(.a(buffered_input), .b(12'b010111101010), .eq(weq1514));
    equaln #(12) e1515(.a(buffered_input), .b(12'b010111101011), .eq(weq1515));
    equaln #(12) e1516(.a(buffered_input), .b(12'b010111101100), .eq(weq1516));
    equaln #(12) e1517(.a(buffered_input), .b(12'b010111101101), .eq(weq1517));
    equaln #(12) e1518(.a(buffered_input), .b(12'b010111101110), .eq(weq1518));
    equaln #(12) e1519(.a(buffered_input), .b(12'b010111101111), .eq(weq1519));
    equaln #(12) e1520(.a(buffered_input), .b(12'b010111110000), .eq(weq1520));
    equaln #(12) e1521(.a(buffered_input), .b(12'b010111110001), .eq(weq1521));
    equaln #(12) e1522(.a(buffered_input), .b(12'b010111110010), .eq(weq1522));
    equaln #(12) e1523(.a(buffered_input), .b(12'b010111110011), .eq(weq1523));
    equaln #(12) e1524(.a(buffered_input), .b(12'b010111110100), .eq(weq1524));
    equaln #(12) e1525(.a(buffered_input), .b(12'b010111110101), .eq(weq1525));
    equaln #(12) e1526(.a(buffered_input), .b(12'b010111110110), .eq(weq1526));
    equaln #(12) e1527(.a(buffered_input), .b(12'b010111110111), .eq(weq1527));
    equaln #(12) e1528(.a(buffered_input), .b(12'b010111111000), .eq(weq1528));
    equaln #(12) e1529(.a(buffered_input), .b(12'b010111111001), .eq(weq1529));
    equaln #(12) e1530(.a(buffered_input), .b(12'b010111111010), .eq(weq1530));
    equaln #(12) e1531(.a(buffered_input), .b(12'b010111111011), .eq(weq1531));
    equaln #(12) e1532(.a(buffered_input), .b(12'b010111111100), .eq(weq1532));
    equaln #(12) e1533(.a(buffered_input), .b(12'b010111111101), .eq(weq1533));
    equaln #(12) e1534(.a(buffered_input), .b(12'b010111111110), .eq(weq1534));
    equaln #(12) e1535(.a(buffered_input), .b(12'b010111111111), .eq(weq1535));
    equaln #(12) e1536(.a(buffered_input), .b(12'b011000000000), .eq(weq1536));
    equaln #(12) e1537(.a(buffered_input), .b(12'b011000000001), .eq(weq1537));
    equaln #(12) e1538(.a(buffered_input), .b(12'b011000000010), .eq(weq1538));
    equaln #(12) e1539(.a(buffered_input), .b(12'b011000000011), .eq(weq1539));
    equaln #(12) e1540(.a(buffered_input), .b(12'b011000000100), .eq(weq1540));
    equaln #(12) e1541(.a(buffered_input), .b(12'b011000000101), .eq(weq1541));
    equaln #(12) e1542(.a(buffered_input), .b(12'b011000000110), .eq(weq1542));
    equaln #(12) e1543(.a(buffered_input), .b(12'b011000000111), .eq(weq1543));
    equaln #(12) e1544(.a(buffered_input), .b(12'b011000001000), .eq(weq1544));
    equaln #(12) e1545(.a(buffered_input), .b(12'b011000001001), .eq(weq1545));
    equaln #(12) e1546(.a(buffered_input), .b(12'b011000001010), .eq(weq1546));
    equaln #(12) e1547(.a(buffered_input), .b(12'b011000001011), .eq(weq1547));
    equaln #(12) e1548(.a(buffered_input), .b(12'b011000001100), .eq(weq1548));
    equaln #(12) e1549(.a(buffered_input), .b(12'b011000001101), .eq(weq1549));
    equaln #(12) e1550(.a(buffered_input), .b(12'b011000001110), .eq(weq1550));
    equaln #(12) e1551(.a(buffered_input), .b(12'b011000001111), .eq(weq1551));
    equaln #(12) e1552(.a(buffered_input), .b(12'b011000010000), .eq(weq1552));
    equaln #(12) e1553(.a(buffered_input), .b(12'b011000010001), .eq(weq1553));
    equaln #(12) e1554(.a(buffered_input), .b(12'b011000010010), .eq(weq1554));
    equaln #(12) e1555(.a(buffered_input), .b(12'b011000010011), .eq(weq1555));
    equaln #(12) e1556(.a(buffered_input), .b(12'b011000010100), .eq(weq1556));
    equaln #(12) e1557(.a(buffered_input), .b(12'b011000010101), .eq(weq1557));
    equaln #(12) e1558(.a(buffered_input), .b(12'b011000010110), .eq(weq1558));
    equaln #(12) e1559(.a(buffered_input), .b(12'b011000010111), .eq(weq1559));
    equaln #(12) e1560(.a(buffered_input), .b(12'b011000011000), .eq(weq1560));
    equaln #(12) e1561(.a(buffered_input), .b(12'b011000011001), .eq(weq1561));
    equaln #(12) e1562(.a(buffered_input), .b(12'b011000011010), .eq(weq1562));
    equaln #(12) e1563(.a(buffered_input), .b(12'b011000011011), .eq(weq1563));
    equaln #(12) e1564(.a(buffered_input), .b(12'b011000011100), .eq(weq1564));
    equaln #(12) e1565(.a(buffered_input), .b(12'b011000011101), .eq(weq1565));
    equaln #(12) e1566(.a(buffered_input), .b(12'b011000011110), .eq(weq1566));
    equaln #(12) e1567(.a(buffered_input), .b(12'b011000011111), .eq(weq1567));
    equaln #(12) e1568(.a(buffered_input), .b(12'b011000100000), .eq(weq1568));
    equaln #(12) e1569(.a(buffered_input), .b(12'b011000100001), .eq(weq1569));
    equaln #(12) e1570(.a(buffered_input), .b(12'b011000100010), .eq(weq1570));
    equaln #(12) e1571(.a(buffered_input), .b(12'b011000100011), .eq(weq1571));
    equaln #(12) e1572(.a(buffered_input), .b(12'b011000100100), .eq(weq1572));
    equaln #(12) e1573(.a(buffered_input), .b(12'b011000100101), .eq(weq1573));
    equaln #(12) e1574(.a(buffered_input), .b(12'b011000100110), .eq(weq1574));
    equaln #(12) e1575(.a(buffered_input), .b(12'b011000100111), .eq(weq1575));
    equaln #(12) e1576(.a(buffered_input), .b(12'b011000101000), .eq(weq1576));
    equaln #(12) e1577(.a(buffered_input), .b(12'b011000101001), .eq(weq1577));
    equaln #(12) e1578(.a(buffered_input), .b(12'b011000101010), .eq(weq1578));
    equaln #(12) e1579(.a(buffered_input), .b(12'b011000101011), .eq(weq1579));
    equaln #(12) e1580(.a(buffered_input), .b(12'b011000101100), .eq(weq1580));
    equaln #(12) e1581(.a(buffered_input), .b(12'b011000101101), .eq(weq1581));
    equaln #(12) e1582(.a(buffered_input), .b(12'b011000101110), .eq(weq1582));
    equaln #(12) e1583(.a(buffered_input), .b(12'b011000101111), .eq(weq1583));
    equaln #(12) e1584(.a(buffered_input), .b(12'b011000110000), .eq(weq1584));
    equaln #(12) e1585(.a(buffered_input), .b(12'b011000110001), .eq(weq1585));
    equaln #(12) e1586(.a(buffered_input), .b(12'b011000110010), .eq(weq1586));
    equaln #(12) e1587(.a(buffered_input), .b(12'b011000110011), .eq(weq1587));
    equaln #(12) e1588(.a(buffered_input), .b(12'b011000110100), .eq(weq1588));
    equaln #(12) e1589(.a(buffered_input), .b(12'b011000110101), .eq(weq1589));
    equaln #(12) e1590(.a(buffered_input), .b(12'b011000110110), .eq(weq1590));
    equaln #(12) e1591(.a(buffered_input), .b(12'b011000110111), .eq(weq1591));
    equaln #(12) e1592(.a(buffered_input), .b(12'b011000111000), .eq(weq1592));
    equaln #(12) e1593(.a(buffered_input), .b(12'b011000111001), .eq(weq1593));
    equaln #(12) e1594(.a(buffered_input), .b(12'b011000111010), .eq(weq1594));
    equaln #(12) e1595(.a(buffered_input), .b(12'b011000111011), .eq(weq1595));
    equaln #(12) e1596(.a(buffered_input), .b(12'b011000111100), .eq(weq1596));
    equaln #(12) e1597(.a(buffered_input), .b(12'b011000111101), .eq(weq1597));
    equaln #(12) e1598(.a(buffered_input), .b(12'b011000111110), .eq(weq1598));
    equaln #(12) e1599(.a(buffered_input), .b(12'b011000111111), .eq(weq1599));
    equaln #(12) e1600(.a(buffered_input), .b(12'b011001000000), .eq(weq1600));
    equaln #(12) e1601(.a(buffered_input), .b(12'b011001000001), .eq(weq1601));
    equaln #(12) e1602(.a(buffered_input), .b(12'b011001000010), .eq(weq1602));
    equaln #(12) e1603(.a(buffered_input), .b(12'b011001000011), .eq(weq1603));
    equaln #(12) e1604(.a(buffered_input), .b(12'b011001000100), .eq(weq1604));
    equaln #(12) e1605(.a(buffered_input), .b(12'b011001000101), .eq(weq1605));
    equaln #(12) e1606(.a(buffered_input), .b(12'b011001000110), .eq(weq1606));
    equaln #(12) e1607(.a(buffered_input), .b(12'b011001000111), .eq(weq1607));
    equaln #(12) e1608(.a(buffered_input), .b(12'b011001001000), .eq(weq1608));
    equaln #(12) e1609(.a(buffered_input), .b(12'b011001001001), .eq(weq1609));
    equaln #(12) e1610(.a(buffered_input), .b(12'b011001001010), .eq(weq1610));
    equaln #(12) e1611(.a(buffered_input), .b(12'b011001001011), .eq(weq1611));
    equaln #(12) e1612(.a(buffered_input), .b(12'b011001001100), .eq(weq1612));
    equaln #(12) e1613(.a(buffered_input), .b(12'b011001001101), .eq(weq1613));
    equaln #(12) e1614(.a(buffered_input), .b(12'b011001001110), .eq(weq1614));
    equaln #(12) e1615(.a(buffered_input), .b(12'b011001001111), .eq(weq1615));
    equaln #(12) e1616(.a(buffered_input), .b(12'b011001010000), .eq(weq1616));
    equaln #(12) e1617(.a(buffered_input), .b(12'b011001010001), .eq(weq1617));
    equaln #(12) e1618(.a(buffered_input), .b(12'b011001010010), .eq(weq1618));
    equaln #(12) e1619(.a(buffered_input), .b(12'b011001010011), .eq(weq1619));
    equaln #(12) e1620(.a(buffered_input), .b(12'b011001010100), .eq(weq1620));
    equaln #(12) e1621(.a(buffered_input), .b(12'b011001010101), .eq(weq1621));
    equaln #(12) e1622(.a(buffered_input), .b(12'b011001010110), .eq(weq1622));
    equaln #(12) e1623(.a(buffered_input), .b(12'b011001010111), .eq(weq1623));
    equaln #(12) e1624(.a(buffered_input), .b(12'b011001011000), .eq(weq1624));
    equaln #(12) e1625(.a(buffered_input), .b(12'b011001011001), .eq(weq1625));
    equaln #(12) e1626(.a(buffered_input), .b(12'b011001011010), .eq(weq1626));
    equaln #(12) e1627(.a(buffered_input), .b(12'b011001011011), .eq(weq1627));
    equaln #(12) e1628(.a(buffered_input), .b(12'b011001011100), .eq(weq1628));
    equaln #(12) e1629(.a(buffered_input), .b(12'b011001011101), .eq(weq1629));
    equaln #(12) e1630(.a(buffered_input), .b(12'b011001011110), .eq(weq1630));
    equaln #(12) e1631(.a(buffered_input), .b(12'b011001011111), .eq(weq1631));
    equaln #(12) e1632(.a(buffered_input), .b(12'b011001100000), .eq(weq1632));
    equaln #(12) e1633(.a(buffered_input), .b(12'b011001100001), .eq(weq1633));
    equaln #(12) e1634(.a(buffered_input), .b(12'b011001100010), .eq(weq1634));
    equaln #(12) e1635(.a(buffered_input), .b(12'b011001100011), .eq(weq1635));
    equaln #(12) e1636(.a(buffered_input), .b(12'b011001100100), .eq(weq1636));
    equaln #(12) e1637(.a(buffered_input), .b(12'b011001100101), .eq(weq1637));
    equaln #(12) e1638(.a(buffered_input), .b(12'b011001100110), .eq(weq1638));
    equaln #(12) e1639(.a(buffered_input), .b(12'b011001100111), .eq(weq1639));
    equaln #(12) e1640(.a(buffered_input), .b(12'b011001101000), .eq(weq1640));
    equaln #(12) e1641(.a(buffered_input), .b(12'b011001101001), .eq(weq1641));
    equaln #(12) e1642(.a(buffered_input), .b(12'b011001101010), .eq(weq1642));
    equaln #(12) e1643(.a(buffered_input), .b(12'b011001101011), .eq(weq1643));
    equaln #(12) e1644(.a(buffered_input), .b(12'b011001101100), .eq(weq1644));
    equaln #(12) e1645(.a(buffered_input), .b(12'b011001101101), .eq(weq1645));
    equaln #(12) e1646(.a(buffered_input), .b(12'b011001101110), .eq(weq1646));
    equaln #(12) e1647(.a(buffered_input), .b(12'b011001101111), .eq(weq1647));
    equaln #(12) e1648(.a(buffered_input), .b(12'b011001110000), .eq(weq1648));
    equaln #(12) e1649(.a(buffered_input), .b(12'b011001110001), .eq(weq1649));
    equaln #(12) e1650(.a(buffered_input), .b(12'b011001110010), .eq(weq1650));
    equaln #(12) e1651(.a(buffered_input), .b(12'b011001110011), .eq(weq1651));
    equaln #(12) e1652(.a(buffered_input), .b(12'b011001110100), .eq(weq1652));
    equaln #(12) e1653(.a(buffered_input), .b(12'b011001110101), .eq(weq1653));
    equaln #(12) e1654(.a(buffered_input), .b(12'b011001110110), .eq(weq1654));
    equaln #(12) e1655(.a(buffered_input), .b(12'b011001110111), .eq(weq1655));
    equaln #(12) e1656(.a(buffered_input), .b(12'b011001111000), .eq(weq1656));
    equaln #(12) e1657(.a(buffered_input), .b(12'b011001111001), .eq(weq1657));
    equaln #(12) e1658(.a(buffered_input), .b(12'b011001111010), .eq(weq1658));
    equaln #(12) e1659(.a(buffered_input), .b(12'b011001111011), .eq(weq1659));
    equaln #(12) e1660(.a(buffered_input), .b(12'b011001111100), .eq(weq1660));
    equaln #(12) e1661(.a(buffered_input), .b(12'b011001111101), .eq(weq1661));
    equaln #(12) e1662(.a(buffered_input), .b(12'b011001111110), .eq(weq1662));
    equaln #(12) e1663(.a(buffered_input), .b(12'b011001111111), .eq(weq1663));
    equaln #(12) e1664(.a(buffered_input), .b(12'b011010000000), .eq(weq1664));
    equaln #(12) e1665(.a(buffered_input), .b(12'b011010000001), .eq(weq1665));
    equaln #(12) e1666(.a(buffered_input), .b(12'b011010000010), .eq(weq1666));
    equaln #(12) e1667(.a(buffered_input), .b(12'b011010000011), .eq(weq1667));
    equaln #(12) e1668(.a(buffered_input), .b(12'b011010000100), .eq(weq1668));
    equaln #(12) e1669(.a(buffered_input), .b(12'b011010000101), .eq(weq1669));
    equaln #(12) e1670(.a(buffered_input), .b(12'b011010000110), .eq(weq1670));
    equaln #(12) e1671(.a(buffered_input), .b(12'b011010000111), .eq(weq1671));
    equaln #(12) e1672(.a(buffered_input), .b(12'b011010001000), .eq(weq1672));
    equaln #(12) e1673(.a(buffered_input), .b(12'b011010001001), .eq(weq1673));
    equaln #(12) e1674(.a(buffered_input), .b(12'b011010001010), .eq(weq1674));
    equaln #(12) e1675(.a(buffered_input), .b(12'b011010001011), .eq(weq1675));
    equaln #(12) e1676(.a(buffered_input), .b(12'b011010001100), .eq(weq1676));
    equaln #(12) e1677(.a(buffered_input), .b(12'b011010001101), .eq(weq1677));
    equaln #(12) e1678(.a(buffered_input), .b(12'b011010001110), .eq(weq1678));
    equaln #(12) e1679(.a(buffered_input), .b(12'b011010001111), .eq(weq1679));
    equaln #(12) e1680(.a(buffered_input), .b(12'b011010010000), .eq(weq1680));
    equaln #(12) e1681(.a(buffered_input), .b(12'b011010010001), .eq(weq1681));
    equaln #(12) e1682(.a(buffered_input), .b(12'b011010010010), .eq(weq1682));
    equaln #(12) e1683(.a(buffered_input), .b(12'b011010010011), .eq(weq1683));
    equaln #(12) e1684(.a(buffered_input), .b(12'b011010010100), .eq(weq1684));
    equaln #(12) e1685(.a(buffered_input), .b(12'b011010010101), .eq(weq1685));
    equaln #(12) e1686(.a(buffered_input), .b(12'b011010010110), .eq(weq1686));
    equaln #(12) e1687(.a(buffered_input), .b(12'b011010010111), .eq(weq1687));
    equaln #(12) e1688(.a(buffered_input), .b(12'b011010011000), .eq(weq1688));
    equaln #(12) e1689(.a(buffered_input), .b(12'b011010011001), .eq(weq1689));
    equaln #(12) e1690(.a(buffered_input), .b(12'b011010011010), .eq(weq1690));
    equaln #(12) e1691(.a(buffered_input), .b(12'b011010011011), .eq(weq1691));
    equaln #(12) e1692(.a(buffered_input), .b(12'b011010011100), .eq(weq1692));
    equaln #(12) e1693(.a(buffered_input), .b(12'b011010011101), .eq(weq1693));
    equaln #(12) e1694(.a(buffered_input), .b(12'b011010011110), .eq(weq1694));
    equaln #(12) e1695(.a(buffered_input), .b(12'b011010011111), .eq(weq1695));
    equaln #(12) e1696(.a(buffered_input), .b(12'b011010100000), .eq(weq1696));
    equaln #(12) e1697(.a(buffered_input), .b(12'b011010100001), .eq(weq1697));
    equaln #(12) e1698(.a(buffered_input), .b(12'b011010100010), .eq(weq1698));
    equaln #(12) e1699(.a(buffered_input), .b(12'b011010100011), .eq(weq1699));
    equaln #(12) e1700(.a(buffered_input), .b(12'b011010100100), .eq(weq1700));
    equaln #(12) e1701(.a(buffered_input), .b(12'b011010100101), .eq(weq1701));
    equaln #(12) e1702(.a(buffered_input), .b(12'b011010100110), .eq(weq1702));
    equaln #(12) e1703(.a(buffered_input), .b(12'b011010100111), .eq(weq1703));
    equaln #(12) e1704(.a(buffered_input), .b(12'b011010101000), .eq(weq1704));
    equaln #(12) e1705(.a(buffered_input), .b(12'b011010101001), .eq(weq1705));
    equaln #(12) e1706(.a(buffered_input), .b(12'b011010101010), .eq(weq1706));
    equaln #(12) e1707(.a(buffered_input), .b(12'b011010101011), .eq(weq1707));
    equaln #(12) e1708(.a(buffered_input), .b(12'b011010101100), .eq(weq1708));
    equaln #(12) e1709(.a(buffered_input), .b(12'b011010101101), .eq(weq1709));
    equaln #(12) e1710(.a(buffered_input), .b(12'b011010101110), .eq(weq1710));
    equaln #(12) e1711(.a(buffered_input), .b(12'b011010101111), .eq(weq1711));
    equaln #(12) e1712(.a(buffered_input), .b(12'b011010110000), .eq(weq1712));
    equaln #(12) e1713(.a(buffered_input), .b(12'b011010110001), .eq(weq1713));
    equaln #(12) e1714(.a(buffered_input), .b(12'b011010110010), .eq(weq1714));
    equaln #(12) e1715(.a(buffered_input), .b(12'b011010110011), .eq(weq1715));
    equaln #(12) e1716(.a(buffered_input), .b(12'b011010110100), .eq(weq1716));
    equaln #(12) e1717(.a(buffered_input), .b(12'b011010110101), .eq(weq1717));
    equaln #(12) e1718(.a(buffered_input), .b(12'b011010110110), .eq(weq1718));
    equaln #(12) e1719(.a(buffered_input), .b(12'b011010110111), .eq(weq1719));
    equaln #(12) e1720(.a(buffered_input), .b(12'b011010111000), .eq(weq1720));
    equaln #(12) e1721(.a(buffered_input), .b(12'b011010111001), .eq(weq1721));
    equaln #(12) e1722(.a(buffered_input), .b(12'b011010111010), .eq(weq1722));
    equaln #(12) e1723(.a(buffered_input), .b(12'b011010111011), .eq(weq1723));
    equaln #(12) e1724(.a(buffered_input), .b(12'b011010111100), .eq(weq1724));
    equaln #(12) e1725(.a(buffered_input), .b(12'b011010111101), .eq(weq1725));
    equaln #(12) e1726(.a(buffered_input), .b(12'b011010111110), .eq(weq1726));
    equaln #(12) e1727(.a(buffered_input), .b(12'b011010111111), .eq(weq1727));
    equaln #(12) e1728(.a(buffered_input), .b(12'b011011000000), .eq(weq1728));
    equaln #(12) e1729(.a(buffered_input), .b(12'b011011000001), .eq(weq1729));
    equaln #(12) e1730(.a(buffered_input), .b(12'b011011000010), .eq(weq1730));
    equaln #(12) e1731(.a(buffered_input), .b(12'b011011000011), .eq(weq1731));
    equaln #(12) e1732(.a(buffered_input), .b(12'b011011000100), .eq(weq1732));
    equaln #(12) e1733(.a(buffered_input), .b(12'b011011000101), .eq(weq1733));
    equaln #(12) e1734(.a(buffered_input), .b(12'b011011000110), .eq(weq1734));
    equaln #(12) e1735(.a(buffered_input), .b(12'b011011000111), .eq(weq1735));
    equaln #(12) e1736(.a(buffered_input), .b(12'b011011001000), .eq(weq1736));
    equaln #(12) e1737(.a(buffered_input), .b(12'b011011001001), .eq(weq1737));
    equaln #(12) e1738(.a(buffered_input), .b(12'b011011001010), .eq(weq1738));
    equaln #(12) e1739(.a(buffered_input), .b(12'b011011001011), .eq(weq1739));
    equaln #(12) e1740(.a(buffered_input), .b(12'b011011001100), .eq(weq1740));
    equaln #(12) e1741(.a(buffered_input), .b(12'b011011001101), .eq(weq1741));
    equaln #(12) e1742(.a(buffered_input), .b(12'b011011001110), .eq(weq1742));
    equaln #(12) e1743(.a(buffered_input), .b(12'b011011001111), .eq(weq1743));
    equaln #(12) e1744(.a(buffered_input), .b(12'b011011010000), .eq(weq1744));
    equaln #(12) e1745(.a(buffered_input), .b(12'b011011010001), .eq(weq1745));
    equaln #(12) e1746(.a(buffered_input), .b(12'b011011010010), .eq(weq1746));
    equaln #(12) e1747(.a(buffered_input), .b(12'b011011010011), .eq(weq1747));
    equaln #(12) e1748(.a(buffered_input), .b(12'b011011010100), .eq(weq1748));
    equaln #(12) e1749(.a(buffered_input), .b(12'b011011010101), .eq(weq1749));
    equaln #(12) e1750(.a(buffered_input), .b(12'b011011010110), .eq(weq1750));
    equaln #(12) e1751(.a(buffered_input), .b(12'b011011010111), .eq(weq1751));
    equaln #(12) e1752(.a(buffered_input), .b(12'b011011011000), .eq(weq1752));
    equaln #(12) e1753(.a(buffered_input), .b(12'b011011011001), .eq(weq1753));
    equaln #(12) e1754(.a(buffered_input), .b(12'b011011011010), .eq(weq1754));
    equaln #(12) e1755(.a(buffered_input), .b(12'b011011011011), .eq(weq1755));
    equaln #(12) e1756(.a(buffered_input), .b(12'b011011011100), .eq(weq1756));
    equaln #(12) e1757(.a(buffered_input), .b(12'b011011011101), .eq(weq1757));
    equaln #(12) e1758(.a(buffered_input), .b(12'b011011011110), .eq(weq1758));
    equaln #(12) e1759(.a(buffered_input), .b(12'b011011011111), .eq(weq1759));
    equaln #(12) e1760(.a(buffered_input), .b(12'b011011100000), .eq(weq1760));
    equaln #(12) e1761(.a(buffered_input), .b(12'b011011100001), .eq(weq1761));
    equaln #(12) e1762(.a(buffered_input), .b(12'b011011100010), .eq(weq1762));
    equaln #(12) e1763(.a(buffered_input), .b(12'b011011100011), .eq(weq1763));
    equaln #(12) e1764(.a(buffered_input), .b(12'b011011100100), .eq(weq1764));
    equaln #(12) e1765(.a(buffered_input), .b(12'b011011100101), .eq(weq1765));
    equaln #(12) e1766(.a(buffered_input), .b(12'b011011100110), .eq(weq1766));
    equaln #(12) e1767(.a(buffered_input), .b(12'b011011100111), .eq(weq1767));
    equaln #(12) e1768(.a(buffered_input), .b(12'b011011101000), .eq(weq1768));
    equaln #(12) e1769(.a(buffered_input), .b(12'b011011101001), .eq(weq1769));
    equaln #(12) e1770(.a(buffered_input), .b(12'b011011101010), .eq(weq1770));
    equaln #(12) e1771(.a(buffered_input), .b(12'b011011101011), .eq(weq1771));
    equaln #(12) e1772(.a(buffered_input), .b(12'b011011101100), .eq(weq1772));
    equaln #(12) e1773(.a(buffered_input), .b(12'b011011101101), .eq(weq1773));
    equaln #(12) e1774(.a(buffered_input), .b(12'b011011101110), .eq(weq1774));
    equaln #(12) e1775(.a(buffered_input), .b(12'b011011101111), .eq(weq1775));
    equaln #(12) e1776(.a(buffered_input), .b(12'b011011110000), .eq(weq1776));
    equaln #(12) e1777(.a(buffered_input), .b(12'b011011110001), .eq(weq1777));
    equaln #(12) e1778(.a(buffered_input), .b(12'b011011110010), .eq(weq1778));
    equaln #(12) e1779(.a(buffered_input), .b(12'b011011110011), .eq(weq1779));
    equaln #(12) e1780(.a(buffered_input), .b(12'b011011110100), .eq(weq1780));
    equaln #(12) e1781(.a(buffered_input), .b(12'b011011110101), .eq(weq1781));
    equaln #(12) e1782(.a(buffered_input), .b(12'b011011110110), .eq(weq1782));
    equaln #(12) e1783(.a(buffered_input), .b(12'b011011110111), .eq(weq1783));
    equaln #(12) e1784(.a(buffered_input), .b(12'b011011111000), .eq(weq1784));
    equaln #(12) e1785(.a(buffered_input), .b(12'b011011111001), .eq(weq1785));
    equaln #(12) e1786(.a(buffered_input), .b(12'b011011111010), .eq(weq1786));
    equaln #(12) e1787(.a(buffered_input), .b(12'b011011111011), .eq(weq1787));
    equaln #(12) e1788(.a(buffered_input), .b(12'b011011111100), .eq(weq1788));
    equaln #(12) e1789(.a(buffered_input), .b(12'b011011111101), .eq(weq1789));
    equaln #(12) e1790(.a(buffered_input), .b(12'b011011111110), .eq(weq1790));
    equaln #(12) e1791(.a(buffered_input), .b(12'b011011111111), .eq(weq1791));
    equaln #(12) e1792(.a(buffered_input), .b(12'b011100000000), .eq(weq1792));
    equaln #(12) e1793(.a(buffered_input), .b(12'b011100000001), .eq(weq1793));
    equaln #(12) e1794(.a(buffered_input), .b(12'b011100000010), .eq(weq1794));
    equaln #(12) e1795(.a(buffered_input), .b(12'b011100000011), .eq(weq1795));
    equaln #(12) e1796(.a(buffered_input), .b(12'b011100000100), .eq(weq1796));
    equaln #(12) e1797(.a(buffered_input), .b(12'b011100000101), .eq(weq1797));
    equaln #(12) e1798(.a(buffered_input), .b(12'b011100000110), .eq(weq1798));
    equaln #(12) e1799(.a(buffered_input), .b(12'b011100000111), .eq(weq1799));
    equaln #(12) e1800(.a(buffered_input), .b(12'b011100001000), .eq(weq1800));
    equaln #(12) e1801(.a(buffered_input), .b(12'b011100001001), .eq(weq1801));
    equaln #(12) e1802(.a(buffered_input), .b(12'b011100001010), .eq(weq1802));
    equaln #(12) e1803(.a(buffered_input), .b(12'b011100001011), .eq(weq1803));
    equaln #(12) e1804(.a(buffered_input), .b(12'b011100001100), .eq(weq1804));
    equaln #(12) e1805(.a(buffered_input), .b(12'b011100001101), .eq(weq1805));
    equaln #(12) e1806(.a(buffered_input), .b(12'b011100001110), .eq(weq1806));
    equaln #(12) e1807(.a(buffered_input), .b(12'b011100001111), .eq(weq1807));
    equaln #(12) e1808(.a(buffered_input), .b(12'b011100010000), .eq(weq1808));
    equaln #(12) e1809(.a(buffered_input), .b(12'b011100010001), .eq(weq1809));
    equaln #(12) e1810(.a(buffered_input), .b(12'b011100010010), .eq(weq1810));
    equaln #(12) e1811(.a(buffered_input), .b(12'b011100010011), .eq(weq1811));
    equaln #(12) e1812(.a(buffered_input), .b(12'b011100010100), .eq(weq1812));
    equaln #(12) e1813(.a(buffered_input), .b(12'b011100010101), .eq(weq1813));
    equaln #(12) e1814(.a(buffered_input), .b(12'b011100010110), .eq(weq1814));
    equaln #(12) e1815(.a(buffered_input), .b(12'b011100010111), .eq(weq1815));
    equaln #(12) e1816(.a(buffered_input), .b(12'b011100011000), .eq(weq1816));
    equaln #(12) e1817(.a(buffered_input), .b(12'b011100011001), .eq(weq1817));
    equaln #(12) e1818(.a(buffered_input), .b(12'b011100011010), .eq(weq1818));
    equaln #(12) e1819(.a(buffered_input), .b(12'b011100011011), .eq(weq1819));
    equaln #(12) e1820(.a(buffered_input), .b(12'b011100011100), .eq(weq1820));
    equaln #(12) e1821(.a(buffered_input), .b(12'b011100011101), .eq(weq1821));
    equaln #(12) e1822(.a(buffered_input), .b(12'b011100011110), .eq(weq1822));
    equaln #(12) e1823(.a(buffered_input), .b(12'b011100011111), .eq(weq1823));
    equaln #(12) e1824(.a(buffered_input), .b(12'b011100100000), .eq(weq1824));
    equaln #(12) e1825(.a(buffered_input), .b(12'b011100100001), .eq(weq1825));
    equaln #(12) e1826(.a(buffered_input), .b(12'b011100100010), .eq(weq1826));
    equaln #(12) e1827(.a(buffered_input), .b(12'b011100100011), .eq(weq1827));
    equaln #(12) e1828(.a(buffered_input), .b(12'b011100100100), .eq(weq1828));
    equaln #(12) e1829(.a(buffered_input), .b(12'b011100100101), .eq(weq1829));
    equaln #(12) e1830(.a(buffered_input), .b(12'b011100100110), .eq(weq1830));
    equaln #(12) e1831(.a(buffered_input), .b(12'b011100100111), .eq(weq1831));
    equaln #(12) e1832(.a(buffered_input), .b(12'b011100101000), .eq(weq1832));
    equaln #(12) e1833(.a(buffered_input), .b(12'b011100101001), .eq(weq1833));
    equaln #(12) e1834(.a(buffered_input), .b(12'b011100101010), .eq(weq1834));
    equaln #(12) e1835(.a(buffered_input), .b(12'b011100101011), .eq(weq1835));
    equaln #(12) e1836(.a(buffered_input), .b(12'b011100101100), .eq(weq1836));
    equaln #(12) e1837(.a(buffered_input), .b(12'b011100101101), .eq(weq1837));
    equaln #(12) e1838(.a(buffered_input), .b(12'b011100101110), .eq(weq1838));
    equaln #(12) e1839(.a(buffered_input), .b(12'b011100101111), .eq(weq1839));
    equaln #(12) e1840(.a(buffered_input), .b(12'b011100110000), .eq(weq1840));
    equaln #(12) e1841(.a(buffered_input), .b(12'b011100110001), .eq(weq1841));
    equaln #(12) e1842(.a(buffered_input), .b(12'b011100110010), .eq(weq1842));
    equaln #(12) e1843(.a(buffered_input), .b(12'b011100110011), .eq(weq1843));
    equaln #(12) e1844(.a(buffered_input), .b(12'b011100110100), .eq(weq1844));
    equaln #(12) e1845(.a(buffered_input), .b(12'b011100110101), .eq(weq1845));
    equaln #(12) e1846(.a(buffered_input), .b(12'b011100110110), .eq(weq1846));
    equaln #(12) e1847(.a(buffered_input), .b(12'b011100110111), .eq(weq1847));
    equaln #(12) e1848(.a(buffered_input), .b(12'b011100111000), .eq(weq1848));
    equaln #(12) e1849(.a(buffered_input), .b(12'b011100111001), .eq(weq1849));
    equaln #(12) e1850(.a(buffered_input), .b(12'b011100111010), .eq(weq1850));
    equaln #(12) e1851(.a(buffered_input), .b(12'b011100111011), .eq(weq1851));
    equaln #(12) e1852(.a(buffered_input), .b(12'b011100111100), .eq(weq1852));
    equaln #(12) e1853(.a(buffered_input), .b(12'b011100111101), .eq(weq1853));
    equaln #(12) e1854(.a(buffered_input), .b(12'b011100111110), .eq(weq1854));
    equaln #(12) e1855(.a(buffered_input), .b(12'b011100111111), .eq(weq1855));
    equaln #(12) e1856(.a(buffered_input), .b(12'b011101000000), .eq(weq1856));
    equaln #(12) e1857(.a(buffered_input), .b(12'b011101000001), .eq(weq1857));
    equaln #(12) e1858(.a(buffered_input), .b(12'b011101000010), .eq(weq1858));
    equaln #(12) e1859(.a(buffered_input), .b(12'b011101000011), .eq(weq1859));
    equaln #(12) e1860(.a(buffered_input), .b(12'b011101000100), .eq(weq1860));
    equaln #(12) e1861(.a(buffered_input), .b(12'b011101000101), .eq(weq1861));
    equaln #(12) e1862(.a(buffered_input), .b(12'b011101000110), .eq(weq1862));
    equaln #(12) e1863(.a(buffered_input), .b(12'b011101000111), .eq(weq1863));
    equaln #(12) e1864(.a(buffered_input), .b(12'b011101001000), .eq(weq1864));
    equaln #(12) e1865(.a(buffered_input), .b(12'b011101001001), .eq(weq1865));
    equaln #(12) e1866(.a(buffered_input), .b(12'b011101001010), .eq(weq1866));
    equaln #(12) e1867(.a(buffered_input), .b(12'b011101001011), .eq(weq1867));
    equaln #(12) e1868(.a(buffered_input), .b(12'b011101001100), .eq(weq1868));
    equaln #(12) e1869(.a(buffered_input), .b(12'b011101001101), .eq(weq1869));
    equaln #(12) e1870(.a(buffered_input), .b(12'b011101001110), .eq(weq1870));
    equaln #(12) e1871(.a(buffered_input), .b(12'b011101001111), .eq(weq1871));
    equaln #(12) e1872(.a(buffered_input), .b(12'b011101010000), .eq(weq1872));
    equaln #(12) e1873(.a(buffered_input), .b(12'b011101010001), .eq(weq1873));
    equaln #(12) e1874(.a(buffered_input), .b(12'b011101010010), .eq(weq1874));
    equaln #(12) e1875(.a(buffered_input), .b(12'b011101010011), .eq(weq1875));
    equaln #(12) e1876(.a(buffered_input), .b(12'b011101010100), .eq(weq1876));
    equaln #(12) e1877(.a(buffered_input), .b(12'b011101010101), .eq(weq1877));
    equaln #(12) e1878(.a(buffered_input), .b(12'b011101010110), .eq(weq1878));
    equaln #(12) e1879(.a(buffered_input), .b(12'b011101010111), .eq(weq1879));
    equaln #(12) e1880(.a(buffered_input), .b(12'b011101011000), .eq(weq1880));
    equaln #(12) e1881(.a(buffered_input), .b(12'b011101011001), .eq(weq1881));
    equaln #(12) e1882(.a(buffered_input), .b(12'b011101011010), .eq(weq1882));
    equaln #(12) e1883(.a(buffered_input), .b(12'b011101011011), .eq(weq1883));
    equaln #(12) e1884(.a(buffered_input), .b(12'b011101011100), .eq(weq1884));
    equaln #(12) e1885(.a(buffered_input), .b(12'b011101011101), .eq(weq1885));
    equaln #(12) e1886(.a(buffered_input), .b(12'b011101011110), .eq(weq1886));
    equaln #(12) e1887(.a(buffered_input), .b(12'b011101011111), .eq(weq1887));
    equaln #(12) e1888(.a(buffered_input), .b(12'b011101100000), .eq(weq1888));
    equaln #(12) e1889(.a(buffered_input), .b(12'b011101100001), .eq(weq1889));
    equaln #(12) e1890(.a(buffered_input), .b(12'b011101100010), .eq(weq1890));
    equaln #(12) e1891(.a(buffered_input), .b(12'b011101100011), .eq(weq1891));
    equaln #(12) e1892(.a(buffered_input), .b(12'b011101100100), .eq(weq1892));
    equaln #(12) e1893(.a(buffered_input), .b(12'b011101100101), .eq(weq1893));
    equaln #(12) e1894(.a(buffered_input), .b(12'b011101100110), .eq(weq1894));
    equaln #(12) e1895(.a(buffered_input), .b(12'b011101100111), .eq(weq1895));
    equaln #(12) e1896(.a(buffered_input), .b(12'b011101101000), .eq(weq1896));
    equaln #(12) e1897(.a(buffered_input), .b(12'b011101101001), .eq(weq1897));
    equaln #(12) e1898(.a(buffered_input), .b(12'b011101101010), .eq(weq1898));
    equaln #(12) e1899(.a(buffered_input), .b(12'b011101101011), .eq(weq1899));
    equaln #(12) e1900(.a(buffered_input), .b(12'b011101101100), .eq(weq1900));
    equaln #(12) e1901(.a(buffered_input), .b(12'b011101101101), .eq(weq1901));
    equaln #(12) e1902(.a(buffered_input), .b(12'b011101101110), .eq(weq1902));
    equaln #(12) e1903(.a(buffered_input), .b(12'b011101101111), .eq(weq1903));
    equaln #(12) e1904(.a(buffered_input), .b(12'b011101110000), .eq(weq1904));
    equaln #(12) e1905(.a(buffered_input), .b(12'b011101110001), .eq(weq1905));
    equaln #(12) e1906(.a(buffered_input), .b(12'b011101110010), .eq(weq1906));
    equaln #(12) e1907(.a(buffered_input), .b(12'b011101110011), .eq(weq1907));
    equaln #(12) e1908(.a(buffered_input), .b(12'b011101110100), .eq(weq1908));
    equaln #(12) e1909(.a(buffered_input), .b(12'b011101110101), .eq(weq1909));
    equaln #(12) e1910(.a(buffered_input), .b(12'b011101110110), .eq(weq1910));
    equaln #(12) e1911(.a(buffered_input), .b(12'b011101110111), .eq(weq1911));
    equaln #(12) e1912(.a(buffered_input), .b(12'b011101111000), .eq(weq1912));
    equaln #(12) e1913(.a(buffered_input), .b(12'b011101111001), .eq(weq1913));
    equaln #(12) e1914(.a(buffered_input), .b(12'b011101111010), .eq(weq1914));
    equaln #(12) e1915(.a(buffered_input), .b(12'b011101111011), .eq(weq1915));
    equaln #(12) e1916(.a(buffered_input), .b(12'b011101111100), .eq(weq1916));
    equaln #(12) e1917(.a(buffered_input), .b(12'b011101111101), .eq(weq1917));
    equaln #(12) e1918(.a(buffered_input), .b(12'b011101111110), .eq(weq1918));
    equaln #(12) e1919(.a(buffered_input), .b(12'b011101111111), .eq(weq1919));
    equaln #(12) e1920(.a(buffered_input), .b(12'b011110000000), .eq(weq1920));
    equaln #(12) e1921(.a(buffered_input), .b(12'b011110000001), .eq(weq1921));
    equaln #(12) e1922(.a(buffered_input), .b(12'b011110000010), .eq(weq1922));
    equaln #(12) e1923(.a(buffered_input), .b(12'b011110000011), .eq(weq1923));
    equaln #(12) e1924(.a(buffered_input), .b(12'b011110000100), .eq(weq1924));
    equaln #(12) e1925(.a(buffered_input), .b(12'b011110000101), .eq(weq1925));
    equaln #(12) e1926(.a(buffered_input), .b(12'b011110000110), .eq(weq1926));
    equaln #(12) e1927(.a(buffered_input), .b(12'b011110000111), .eq(weq1927));
    equaln #(12) e1928(.a(buffered_input), .b(12'b011110001000), .eq(weq1928));
    equaln #(12) e1929(.a(buffered_input), .b(12'b011110001001), .eq(weq1929));
    equaln #(12) e1930(.a(buffered_input), .b(12'b011110001010), .eq(weq1930));
    equaln #(12) e1931(.a(buffered_input), .b(12'b011110001011), .eq(weq1931));
    equaln #(12) e1932(.a(buffered_input), .b(12'b011110001100), .eq(weq1932));
    equaln #(12) e1933(.a(buffered_input), .b(12'b011110001101), .eq(weq1933));
    equaln #(12) e1934(.a(buffered_input), .b(12'b011110001110), .eq(weq1934));
    equaln #(12) e1935(.a(buffered_input), .b(12'b011110001111), .eq(weq1935));
    equaln #(12) e1936(.a(buffered_input), .b(12'b011110010000), .eq(weq1936));
    equaln #(12) e1937(.a(buffered_input), .b(12'b011110010001), .eq(weq1937));
    equaln #(12) e1938(.a(buffered_input), .b(12'b011110010010), .eq(weq1938));
    equaln #(12) e1939(.a(buffered_input), .b(12'b011110010011), .eq(weq1939));
    equaln #(12) e1940(.a(buffered_input), .b(12'b011110010100), .eq(weq1940));
    equaln #(12) e1941(.a(buffered_input), .b(12'b011110010101), .eq(weq1941));
    equaln #(12) e1942(.a(buffered_input), .b(12'b011110010110), .eq(weq1942));
    equaln #(12) e1943(.a(buffered_input), .b(12'b011110010111), .eq(weq1943));
    equaln #(12) e1944(.a(buffered_input), .b(12'b011110011000), .eq(weq1944));
    equaln #(12) e1945(.a(buffered_input), .b(12'b011110011001), .eq(weq1945));
    equaln #(12) e1946(.a(buffered_input), .b(12'b011110011010), .eq(weq1946));
    equaln #(12) e1947(.a(buffered_input), .b(12'b011110011011), .eq(weq1947));
    equaln #(12) e1948(.a(buffered_input), .b(12'b011110011100), .eq(weq1948));
    equaln #(12) e1949(.a(buffered_input), .b(12'b011110011101), .eq(weq1949));
    equaln #(12) e1950(.a(buffered_input), .b(12'b011110011110), .eq(weq1950));
    equaln #(12) e1951(.a(buffered_input), .b(12'b011110011111), .eq(weq1951));
    equaln #(12) e1952(.a(buffered_input), .b(12'b011110100000), .eq(weq1952));
    equaln #(12) e1953(.a(buffered_input), .b(12'b011110100001), .eq(weq1953));
    equaln #(12) e1954(.a(buffered_input), .b(12'b011110100010), .eq(weq1954));
    equaln #(12) e1955(.a(buffered_input), .b(12'b011110100011), .eq(weq1955));
    equaln #(12) e1956(.a(buffered_input), .b(12'b011110100100), .eq(weq1956));
    equaln #(12) e1957(.a(buffered_input), .b(12'b011110100101), .eq(weq1957));
    equaln #(12) e1958(.a(buffered_input), .b(12'b011110100110), .eq(weq1958));
    equaln #(12) e1959(.a(buffered_input), .b(12'b011110100111), .eq(weq1959));
    equaln #(12) e1960(.a(buffered_input), .b(12'b011110101000), .eq(weq1960));
    equaln #(12) e1961(.a(buffered_input), .b(12'b011110101001), .eq(weq1961));
    equaln #(12) e1962(.a(buffered_input), .b(12'b011110101010), .eq(weq1962));
    equaln #(12) e1963(.a(buffered_input), .b(12'b011110101011), .eq(weq1963));
    equaln #(12) e1964(.a(buffered_input), .b(12'b011110101100), .eq(weq1964));
    equaln #(12) e1965(.a(buffered_input), .b(12'b011110101101), .eq(weq1965));
    equaln #(12) e1966(.a(buffered_input), .b(12'b011110101110), .eq(weq1966));
    equaln #(12) e1967(.a(buffered_input), .b(12'b011110101111), .eq(weq1967));
    equaln #(12) e1968(.a(buffered_input), .b(12'b011110110000), .eq(weq1968));
    equaln #(12) e1969(.a(buffered_input), .b(12'b011110110001), .eq(weq1969));
    equaln #(12) e1970(.a(buffered_input), .b(12'b011110110010), .eq(weq1970));
    equaln #(12) e1971(.a(buffered_input), .b(12'b011110110011), .eq(weq1971));
    equaln #(12) e1972(.a(buffered_input), .b(12'b011110110100), .eq(weq1972));
    equaln #(12) e1973(.a(buffered_input), .b(12'b011110110101), .eq(weq1973));
    equaln #(12) e1974(.a(buffered_input), .b(12'b011110110110), .eq(weq1974));
    equaln #(12) e1975(.a(buffered_input), .b(12'b011110110111), .eq(weq1975));
    equaln #(12) e1976(.a(buffered_input), .b(12'b011110111000), .eq(weq1976));
    equaln #(12) e1977(.a(buffered_input), .b(12'b011110111001), .eq(weq1977));
    equaln #(12) e1978(.a(buffered_input), .b(12'b011110111010), .eq(weq1978));
    equaln #(12) e1979(.a(buffered_input), .b(12'b011110111011), .eq(weq1979));
    equaln #(12) e1980(.a(buffered_input), .b(12'b011110111100), .eq(weq1980));
    equaln #(12) e1981(.a(buffered_input), .b(12'b011110111101), .eq(weq1981));
    equaln #(12) e1982(.a(buffered_input), .b(12'b011110111110), .eq(weq1982));
    equaln #(12) e1983(.a(buffered_input), .b(12'b011110111111), .eq(weq1983));
    equaln #(12) e1984(.a(buffered_input), .b(12'b011111000000), .eq(weq1984));
    equaln #(12) e1985(.a(buffered_input), .b(12'b011111000001), .eq(weq1985));
    equaln #(12) e1986(.a(buffered_input), .b(12'b011111000010), .eq(weq1986));
    equaln #(12) e1987(.a(buffered_input), .b(12'b011111000011), .eq(weq1987));
    equaln #(12) e1988(.a(buffered_input), .b(12'b011111000100), .eq(weq1988));
    equaln #(12) e1989(.a(buffered_input), .b(12'b011111000101), .eq(weq1989));
    equaln #(12) e1990(.a(buffered_input), .b(12'b011111000110), .eq(weq1990));
    equaln #(12) e1991(.a(buffered_input), .b(12'b011111000111), .eq(weq1991));
    equaln #(12) e1992(.a(buffered_input), .b(12'b011111001000), .eq(weq1992));
    equaln #(12) e1993(.a(buffered_input), .b(12'b011111001001), .eq(weq1993));
    equaln #(12) e1994(.a(buffered_input), .b(12'b011111001010), .eq(weq1994));
    equaln #(12) e1995(.a(buffered_input), .b(12'b011111001011), .eq(weq1995));
    equaln #(12) e1996(.a(buffered_input), .b(12'b011111001100), .eq(weq1996));
    equaln #(12) e1997(.a(buffered_input), .b(12'b011111001101), .eq(weq1997));
    equaln #(12) e1998(.a(buffered_input), .b(12'b011111001110), .eq(weq1998));
    equaln #(12) e1999(.a(buffered_input), .b(12'b011111001111), .eq(weq1999));
    equaln #(12) e2000(.a(buffered_input), .b(12'b011111010000), .eq(weq2000));
    equaln #(12) e2001(.a(buffered_input), .b(12'b011111010001), .eq(weq2001));
    equaln #(12) e2002(.a(buffered_input), .b(12'b011111010010), .eq(weq2002));
    equaln #(12) e2003(.a(buffered_input), .b(12'b011111010011), .eq(weq2003));
    equaln #(12) e2004(.a(buffered_input), .b(12'b011111010100), .eq(weq2004));
    equaln #(12) e2005(.a(buffered_input), .b(12'b011111010101), .eq(weq2005));
    equaln #(12) e2006(.a(buffered_input), .b(12'b011111010110), .eq(weq2006));
    equaln #(12) e2007(.a(buffered_input), .b(12'b011111010111), .eq(weq2007));
    equaln #(12) e2008(.a(buffered_input), .b(12'b011111011000), .eq(weq2008));
    equaln #(12) e2009(.a(buffered_input), .b(12'b011111011001), .eq(weq2009));
    equaln #(12) e2010(.a(buffered_input), .b(12'b011111011010), .eq(weq2010));
    equaln #(12) e2011(.a(buffered_input), .b(12'b011111011011), .eq(weq2011));
    equaln #(12) e2012(.a(buffered_input), .b(12'b011111011100), .eq(weq2012));
    equaln #(12) e2013(.a(buffered_input), .b(12'b011111011101), .eq(weq2013));
    equaln #(12) e2014(.a(buffered_input), .b(12'b011111011110), .eq(weq2014));
    equaln #(12) e2015(.a(buffered_input), .b(12'b011111011111), .eq(weq2015));
    equaln #(12) e2016(.a(buffered_input), .b(12'b011111100000), .eq(weq2016));
    equaln #(12) e2017(.a(buffered_input), .b(12'b011111100001), .eq(weq2017));
    equaln #(12) e2018(.a(buffered_input), .b(12'b011111100010), .eq(weq2018));
    equaln #(12) e2019(.a(buffered_input), .b(12'b011111100011), .eq(weq2019));
    equaln #(12) e2020(.a(buffered_input), .b(12'b011111100100), .eq(weq2020));
    equaln #(12) e2021(.a(buffered_input), .b(12'b011111100101), .eq(weq2021));
    equaln #(12) e2022(.a(buffered_input), .b(12'b011111100110), .eq(weq2022));
    equaln #(12) e2023(.a(buffered_input), .b(12'b011111100111), .eq(weq2023));
    equaln #(12) e2024(.a(buffered_input), .b(12'b011111101000), .eq(weq2024));
    equaln #(12) e2025(.a(buffered_input), .b(12'b011111101001), .eq(weq2025));
    equaln #(12) e2026(.a(buffered_input), .b(12'b011111101010), .eq(weq2026));
    equaln #(12) e2027(.a(buffered_input), .b(12'b011111101011), .eq(weq2027));
    equaln #(12) e2028(.a(buffered_input), .b(12'b011111101100), .eq(weq2028));
    equaln #(12) e2029(.a(buffered_input), .b(12'b011111101101), .eq(weq2029));
    equaln #(12) e2030(.a(buffered_input), .b(12'b011111101110), .eq(weq2030));
    equaln #(12) e2031(.a(buffered_input), .b(12'b011111101111), .eq(weq2031));
    equaln #(12) e2032(.a(buffered_input), .b(12'b011111110000), .eq(weq2032));
    equaln #(12) e2033(.a(buffered_input), .b(12'b011111110001), .eq(weq2033));
    equaln #(12) e2034(.a(buffered_input), .b(12'b011111110010), .eq(weq2034));
    equaln #(12) e2035(.a(buffered_input), .b(12'b011111110011), .eq(weq2035));
    equaln #(12) e2036(.a(buffered_input), .b(12'b011111110100), .eq(weq2036));
    equaln #(12) e2037(.a(buffered_input), .b(12'b011111110101), .eq(weq2037));
    equaln #(12) e2038(.a(buffered_input), .b(12'b011111110110), .eq(weq2038));
    equaln #(12) e2039(.a(buffered_input), .b(12'b011111110111), .eq(weq2039));
    equaln #(12) e2040(.a(buffered_input), .b(12'b011111111000), .eq(weq2040));
    equaln #(12) e2041(.a(buffered_input), .b(12'b011111111001), .eq(weq2041));
    equaln #(12) e2042(.a(buffered_input), .b(12'b011111111010), .eq(weq2042));
    equaln #(12) e2043(.a(buffered_input), .b(12'b011111111011), .eq(weq2043));
    equaln #(12) e2044(.a(buffered_input), .b(12'b011111111100), .eq(weq2044));
    equaln #(12) e2045(.a(buffered_input), .b(12'b011111111101), .eq(weq2045));
    equaln #(12) e2046(.a(buffered_input), .b(12'b011111111110), .eq(weq2046));
    equaln #(12) e2047(.a(buffered_input), .b(12'b011111111111), .eq(weq2047));
    equaln #(12) e2048(.a(buffered_input), .b(12'b100000000000), .eq(weq2048));
    equaln #(12) e2049(.a(buffered_input), .b(12'b100000000001), .eq(weq2049));
    equaln #(12) e2050(.a(buffered_input), .b(12'b100000000010), .eq(weq2050));
    equaln #(12) e2051(.a(buffered_input), .b(12'b100000000011), .eq(weq2051));
    equaln #(12) e2052(.a(buffered_input), .b(12'b100000000100), .eq(weq2052));
    equaln #(12) e2053(.a(buffered_input), .b(12'b100000000101), .eq(weq2053));
    equaln #(12) e2054(.a(buffered_input), .b(12'b100000000110), .eq(weq2054));
    equaln #(12) e2055(.a(buffered_input), .b(12'b100000000111), .eq(weq2055));
    equaln #(12) e2056(.a(buffered_input), .b(12'b100000001000), .eq(weq2056));
    equaln #(12) e2057(.a(buffered_input), .b(12'b100000001001), .eq(weq2057));
    equaln #(12) e2058(.a(buffered_input), .b(12'b100000001010), .eq(weq2058));
    equaln #(12) e2059(.a(buffered_input), .b(12'b100000001011), .eq(weq2059));
    equaln #(12) e2060(.a(buffered_input), .b(12'b100000001100), .eq(weq2060));
    equaln #(12) e2061(.a(buffered_input), .b(12'b100000001101), .eq(weq2061));
    equaln #(12) e2062(.a(buffered_input), .b(12'b100000001110), .eq(weq2062));
    equaln #(12) e2063(.a(buffered_input), .b(12'b100000001111), .eq(weq2063));
    equaln #(12) e2064(.a(buffered_input), .b(12'b100000010000), .eq(weq2064));
    equaln #(12) e2065(.a(buffered_input), .b(12'b100000010001), .eq(weq2065));
    equaln #(12) e2066(.a(buffered_input), .b(12'b100000010010), .eq(weq2066));
    equaln #(12) e2067(.a(buffered_input), .b(12'b100000010011), .eq(weq2067));
    equaln #(12) e2068(.a(buffered_input), .b(12'b100000010100), .eq(weq2068));
    equaln #(12) e2069(.a(buffered_input), .b(12'b100000010101), .eq(weq2069));
    equaln #(12) e2070(.a(buffered_input), .b(12'b100000010110), .eq(weq2070));
    equaln #(12) e2071(.a(buffered_input), .b(12'b100000010111), .eq(weq2071));
    equaln #(12) e2072(.a(buffered_input), .b(12'b100000011000), .eq(weq2072));
    equaln #(12) e2073(.a(buffered_input), .b(12'b100000011001), .eq(weq2073));
    equaln #(12) e2074(.a(buffered_input), .b(12'b100000011010), .eq(weq2074));
    equaln #(12) e2075(.a(buffered_input), .b(12'b100000011011), .eq(weq2075));
    equaln #(12) e2076(.a(buffered_input), .b(12'b100000011100), .eq(weq2076));
    equaln #(12) e2077(.a(buffered_input), .b(12'b100000011101), .eq(weq2077));
    equaln #(12) e2078(.a(buffered_input), .b(12'b100000011110), .eq(weq2078));
    equaln #(12) e2079(.a(buffered_input), .b(12'b100000011111), .eq(weq2079));
    equaln #(12) e2080(.a(buffered_input), .b(12'b100000100000), .eq(weq2080));
    equaln #(12) e2081(.a(buffered_input), .b(12'b100000100001), .eq(weq2081));
    equaln #(12) e2082(.a(buffered_input), .b(12'b100000100010), .eq(weq2082));
    equaln #(12) e2083(.a(buffered_input), .b(12'b100000100011), .eq(weq2083));
    equaln #(12) e2084(.a(buffered_input), .b(12'b100000100100), .eq(weq2084));
    equaln #(12) e2085(.a(buffered_input), .b(12'b100000100101), .eq(weq2085));
    equaln #(12) e2086(.a(buffered_input), .b(12'b100000100110), .eq(weq2086));
    equaln #(12) e2087(.a(buffered_input), .b(12'b100000100111), .eq(weq2087));
    equaln #(12) e2088(.a(buffered_input), .b(12'b100000101000), .eq(weq2088));
    equaln #(12) e2089(.a(buffered_input), .b(12'b100000101001), .eq(weq2089));
    equaln #(12) e2090(.a(buffered_input), .b(12'b100000101010), .eq(weq2090));
    equaln #(12) e2091(.a(buffered_input), .b(12'b100000101011), .eq(weq2091));
    equaln #(12) e2092(.a(buffered_input), .b(12'b100000101100), .eq(weq2092));
    equaln #(12) e2093(.a(buffered_input), .b(12'b100000101101), .eq(weq2093));
    equaln #(12) e2094(.a(buffered_input), .b(12'b100000101110), .eq(weq2094));
    equaln #(12) e2095(.a(buffered_input), .b(12'b100000101111), .eq(weq2095));
    equaln #(12) e2096(.a(buffered_input), .b(12'b100000110000), .eq(weq2096));
    equaln #(12) e2097(.a(buffered_input), .b(12'b100000110001), .eq(weq2097));
    equaln #(12) e2098(.a(buffered_input), .b(12'b100000110010), .eq(weq2098));
    equaln #(12) e2099(.a(buffered_input), .b(12'b100000110011), .eq(weq2099));
    equaln #(12) e2100(.a(buffered_input), .b(12'b100000110100), .eq(weq2100));
    equaln #(12) e2101(.a(buffered_input), .b(12'b100000110101), .eq(weq2101));
    equaln #(12) e2102(.a(buffered_input), .b(12'b100000110110), .eq(weq2102));
    equaln #(12) e2103(.a(buffered_input), .b(12'b100000110111), .eq(weq2103));
    equaln #(12) e2104(.a(buffered_input), .b(12'b100000111000), .eq(weq2104));
    equaln #(12) e2105(.a(buffered_input), .b(12'b100000111001), .eq(weq2105));
    equaln #(12) e2106(.a(buffered_input), .b(12'b100000111010), .eq(weq2106));
    equaln #(12) e2107(.a(buffered_input), .b(12'b100000111011), .eq(weq2107));
    equaln #(12) e2108(.a(buffered_input), .b(12'b100000111100), .eq(weq2108));
    equaln #(12) e2109(.a(buffered_input), .b(12'b100000111101), .eq(weq2109));
    equaln #(12) e2110(.a(buffered_input), .b(12'b100000111110), .eq(weq2110));
    equaln #(12) e2111(.a(buffered_input), .b(12'b100000111111), .eq(weq2111));
    equaln #(12) e2112(.a(buffered_input), .b(12'b100001000000), .eq(weq2112));
    equaln #(12) e2113(.a(buffered_input), .b(12'b100001000001), .eq(weq2113));
    equaln #(12) e2114(.a(buffered_input), .b(12'b100001000010), .eq(weq2114));
    equaln #(12) e2115(.a(buffered_input), .b(12'b100001000011), .eq(weq2115));
    equaln #(12) e2116(.a(buffered_input), .b(12'b100001000100), .eq(weq2116));
    equaln #(12) e2117(.a(buffered_input), .b(12'b100001000101), .eq(weq2117));
    equaln #(12) e2118(.a(buffered_input), .b(12'b100001000110), .eq(weq2118));
    equaln #(12) e2119(.a(buffered_input), .b(12'b100001000111), .eq(weq2119));
    equaln #(12) e2120(.a(buffered_input), .b(12'b100001001000), .eq(weq2120));
    equaln #(12) e2121(.a(buffered_input), .b(12'b100001001001), .eq(weq2121));
    equaln #(12) e2122(.a(buffered_input), .b(12'b100001001010), .eq(weq2122));
    equaln #(12) e2123(.a(buffered_input), .b(12'b100001001011), .eq(weq2123));
    equaln #(12) e2124(.a(buffered_input), .b(12'b100001001100), .eq(weq2124));
    equaln #(12) e2125(.a(buffered_input), .b(12'b100001001101), .eq(weq2125));
    equaln #(12) e2126(.a(buffered_input), .b(12'b100001001110), .eq(weq2126));
    equaln #(12) e2127(.a(buffered_input), .b(12'b100001001111), .eq(weq2127));
    equaln #(12) e2128(.a(buffered_input), .b(12'b100001010000), .eq(weq2128));
    equaln #(12) e2129(.a(buffered_input), .b(12'b100001010001), .eq(weq2129));
    equaln #(12) e2130(.a(buffered_input), .b(12'b100001010010), .eq(weq2130));
    equaln #(12) e2131(.a(buffered_input), .b(12'b100001010011), .eq(weq2131));
    equaln #(12) e2132(.a(buffered_input), .b(12'b100001010100), .eq(weq2132));
    equaln #(12) e2133(.a(buffered_input), .b(12'b100001010101), .eq(weq2133));
    equaln #(12) e2134(.a(buffered_input), .b(12'b100001010110), .eq(weq2134));
    equaln #(12) e2135(.a(buffered_input), .b(12'b100001010111), .eq(weq2135));
    equaln #(12) e2136(.a(buffered_input), .b(12'b100001011000), .eq(weq2136));
    equaln #(12) e2137(.a(buffered_input), .b(12'b100001011001), .eq(weq2137));
    equaln #(12) e2138(.a(buffered_input), .b(12'b100001011010), .eq(weq2138));
    equaln #(12) e2139(.a(buffered_input), .b(12'b100001011011), .eq(weq2139));
    equaln #(12) e2140(.a(buffered_input), .b(12'b100001011100), .eq(weq2140));
    equaln #(12) e2141(.a(buffered_input), .b(12'b100001011101), .eq(weq2141));
    equaln #(12) e2142(.a(buffered_input), .b(12'b100001011110), .eq(weq2142));
    equaln #(12) e2143(.a(buffered_input), .b(12'b100001011111), .eq(weq2143));
    equaln #(12) e2144(.a(buffered_input), .b(12'b100001100000), .eq(weq2144));
    equaln #(12) e2145(.a(buffered_input), .b(12'b100001100001), .eq(weq2145));
    equaln #(12) e2146(.a(buffered_input), .b(12'b100001100010), .eq(weq2146));
    equaln #(12) e2147(.a(buffered_input), .b(12'b100001100011), .eq(weq2147));
    equaln #(12) e2148(.a(buffered_input), .b(12'b100001100100), .eq(weq2148));
    equaln #(12) e2149(.a(buffered_input), .b(12'b100001100101), .eq(weq2149));
    equaln #(12) e2150(.a(buffered_input), .b(12'b100001100110), .eq(weq2150));
    equaln #(12) e2151(.a(buffered_input), .b(12'b100001100111), .eq(weq2151));
    equaln #(12) e2152(.a(buffered_input), .b(12'b100001101000), .eq(weq2152));
    equaln #(12) e2153(.a(buffered_input), .b(12'b100001101001), .eq(weq2153));
    equaln #(12) e2154(.a(buffered_input), .b(12'b100001101010), .eq(weq2154));
    equaln #(12) e2155(.a(buffered_input), .b(12'b100001101011), .eq(weq2155));
    equaln #(12) e2156(.a(buffered_input), .b(12'b100001101100), .eq(weq2156));
    equaln #(12) e2157(.a(buffered_input), .b(12'b100001101101), .eq(weq2157));
    equaln #(12) e2158(.a(buffered_input), .b(12'b100001101110), .eq(weq2158));
    equaln #(12) e2159(.a(buffered_input), .b(12'b100001101111), .eq(weq2159));
    equaln #(12) e2160(.a(buffered_input), .b(12'b100001110000), .eq(weq2160));
    equaln #(12) e2161(.a(buffered_input), .b(12'b100001110001), .eq(weq2161));
    equaln #(12) e2162(.a(buffered_input), .b(12'b100001110010), .eq(weq2162));
    equaln #(12) e2163(.a(buffered_input), .b(12'b100001110011), .eq(weq2163));
    equaln #(12) e2164(.a(buffered_input), .b(12'b100001110100), .eq(weq2164));
    equaln #(12) e2165(.a(buffered_input), .b(12'b100001110101), .eq(weq2165));
    equaln #(12) e2166(.a(buffered_input), .b(12'b100001110110), .eq(weq2166));
    equaln #(12) e2167(.a(buffered_input), .b(12'b100001110111), .eq(weq2167));
    equaln #(12) e2168(.a(buffered_input), .b(12'b100001111000), .eq(weq2168));
    equaln #(12) e2169(.a(buffered_input), .b(12'b100001111001), .eq(weq2169));
    equaln #(12) e2170(.a(buffered_input), .b(12'b100001111010), .eq(weq2170));
    equaln #(12) e2171(.a(buffered_input), .b(12'b100001111011), .eq(weq2171));
    equaln #(12) e2172(.a(buffered_input), .b(12'b100001111100), .eq(weq2172));
    equaln #(12) e2173(.a(buffered_input), .b(12'b100001111101), .eq(weq2173));
    equaln #(12) e2174(.a(buffered_input), .b(12'b100001111110), .eq(weq2174));
    equaln #(12) e2175(.a(buffered_input), .b(12'b100001111111), .eq(weq2175));
    equaln #(12) e2176(.a(buffered_input), .b(12'b100010000000), .eq(weq2176));
    equaln #(12) e2177(.a(buffered_input), .b(12'b100010000001), .eq(weq2177));
    equaln #(12) e2178(.a(buffered_input), .b(12'b100010000010), .eq(weq2178));
    equaln #(12) e2179(.a(buffered_input), .b(12'b100010000011), .eq(weq2179));
    equaln #(12) e2180(.a(buffered_input), .b(12'b100010000100), .eq(weq2180));
    equaln #(12) e2181(.a(buffered_input), .b(12'b100010000101), .eq(weq2181));
    equaln #(12) e2182(.a(buffered_input), .b(12'b100010000110), .eq(weq2182));
    equaln #(12) e2183(.a(buffered_input), .b(12'b100010000111), .eq(weq2183));
    equaln #(12) e2184(.a(buffered_input), .b(12'b100010001000), .eq(weq2184));
    equaln #(12) e2185(.a(buffered_input), .b(12'b100010001001), .eq(weq2185));
    equaln #(12) e2186(.a(buffered_input), .b(12'b100010001010), .eq(weq2186));
    equaln #(12) e2187(.a(buffered_input), .b(12'b100010001011), .eq(weq2187));
    equaln #(12) e2188(.a(buffered_input), .b(12'b100010001100), .eq(weq2188));
    equaln #(12) e2189(.a(buffered_input), .b(12'b100010001101), .eq(weq2189));
    equaln #(12) e2190(.a(buffered_input), .b(12'b100010001110), .eq(weq2190));
    equaln #(12) e2191(.a(buffered_input), .b(12'b100010001111), .eq(weq2191));
    equaln #(12) e2192(.a(buffered_input), .b(12'b100010010000), .eq(weq2192));
    equaln #(12) e2193(.a(buffered_input), .b(12'b100010010001), .eq(weq2193));
    equaln #(12) e2194(.a(buffered_input), .b(12'b100010010010), .eq(weq2194));
    equaln #(12) e2195(.a(buffered_input), .b(12'b100010010011), .eq(weq2195));
    equaln #(12) e2196(.a(buffered_input), .b(12'b100010010100), .eq(weq2196));
    equaln #(12) e2197(.a(buffered_input), .b(12'b100010010101), .eq(weq2197));
    equaln #(12) e2198(.a(buffered_input), .b(12'b100010010110), .eq(weq2198));
    equaln #(12) e2199(.a(buffered_input), .b(12'b100010010111), .eq(weq2199));
    equaln #(12) e2200(.a(buffered_input), .b(12'b100010011000), .eq(weq2200));
    equaln #(12) e2201(.a(buffered_input), .b(12'b100010011001), .eq(weq2201));
    equaln #(12) e2202(.a(buffered_input), .b(12'b100010011010), .eq(weq2202));
    equaln #(12) e2203(.a(buffered_input), .b(12'b100010011011), .eq(weq2203));
    equaln #(12) e2204(.a(buffered_input), .b(12'b100010011100), .eq(weq2204));
    equaln #(12) e2205(.a(buffered_input), .b(12'b100010011101), .eq(weq2205));
    equaln #(12) e2206(.a(buffered_input), .b(12'b100010011110), .eq(weq2206));
    equaln #(12) e2207(.a(buffered_input), .b(12'b100010011111), .eq(weq2207));
    equaln #(12) e2208(.a(buffered_input), .b(12'b100010100000), .eq(weq2208));
    equaln #(12) e2209(.a(buffered_input), .b(12'b100010100001), .eq(weq2209));
    equaln #(12) e2210(.a(buffered_input), .b(12'b100010100010), .eq(weq2210));
    equaln #(12) e2211(.a(buffered_input), .b(12'b100010100011), .eq(weq2211));
    equaln #(12) e2212(.a(buffered_input), .b(12'b100010100100), .eq(weq2212));
    equaln #(12) e2213(.a(buffered_input), .b(12'b100010100101), .eq(weq2213));
    equaln #(12) e2214(.a(buffered_input), .b(12'b100010100110), .eq(weq2214));
    equaln #(12) e2215(.a(buffered_input), .b(12'b100010100111), .eq(weq2215));
    equaln #(12) e2216(.a(buffered_input), .b(12'b100010101000), .eq(weq2216));
    equaln #(12) e2217(.a(buffered_input), .b(12'b100010101001), .eq(weq2217));
    equaln #(12) e2218(.a(buffered_input), .b(12'b100010101010), .eq(weq2218));
    equaln #(12) e2219(.a(buffered_input), .b(12'b100010101011), .eq(weq2219));
    equaln #(12) e2220(.a(buffered_input), .b(12'b100010101100), .eq(weq2220));
    equaln #(12) e2221(.a(buffered_input), .b(12'b100010101101), .eq(weq2221));
    equaln #(12) e2222(.a(buffered_input), .b(12'b100010101110), .eq(weq2222));
    equaln #(12) e2223(.a(buffered_input), .b(12'b100010101111), .eq(weq2223));
    equaln #(12) e2224(.a(buffered_input), .b(12'b100010110000), .eq(weq2224));
    equaln #(12) e2225(.a(buffered_input), .b(12'b100010110001), .eq(weq2225));
    equaln #(12) e2226(.a(buffered_input), .b(12'b100010110010), .eq(weq2226));
    equaln #(12) e2227(.a(buffered_input), .b(12'b100010110011), .eq(weq2227));
    equaln #(12) e2228(.a(buffered_input), .b(12'b100010110100), .eq(weq2228));
    equaln #(12) e2229(.a(buffered_input), .b(12'b100010110101), .eq(weq2229));
    equaln #(12) e2230(.a(buffered_input), .b(12'b100010110110), .eq(weq2230));
    equaln #(12) e2231(.a(buffered_input), .b(12'b100010110111), .eq(weq2231));
    equaln #(12) e2232(.a(buffered_input), .b(12'b100010111000), .eq(weq2232));
    equaln #(12) e2233(.a(buffered_input), .b(12'b100010111001), .eq(weq2233));
    equaln #(12) e2234(.a(buffered_input), .b(12'b100010111010), .eq(weq2234));
    equaln #(12) e2235(.a(buffered_input), .b(12'b100010111011), .eq(weq2235));
    equaln #(12) e2236(.a(buffered_input), .b(12'b100010111100), .eq(weq2236));
    equaln #(12) e2237(.a(buffered_input), .b(12'b100010111101), .eq(weq2237));
    equaln #(12) e2238(.a(buffered_input), .b(12'b100010111110), .eq(weq2238));
    equaln #(12) e2239(.a(buffered_input), .b(12'b100010111111), .eq(weq2239));
    equaln #(12) e2240(.a(buffered_input), .b(12'b100011000000), .eq(weq2240));
    equaln #(12) e2241(.a(buffered_input), .b(12'b100011000001), .eq(weq2241));
    equaln #(12) e2242(.a(buffered_input), .b(12'b100011000010), .eq(weq2242));
    equaln #(12) e2243(.a(buffered_input), .b(12'b100011000011), .eq(weq2243));
    equaln #(12) e2244(.a(buffered_input), .b(12'b100011000100), .eq(weq2244));
    equaln #(12) e2245(.a(buffered_input), .b(12'b100011000101), .eq(weq2245));
    equaln #(12) e2246(.a(buffered_input), .b(12'b100011000110), .eq(weq2246));
    equaln #(12) e2247(.a(buffered_input), .b(12'b100011000111), .eq(weq2247));
    equaln #(12) e2248(.a(buffered_input), .b(12'b100011001000), .eq(weq2248));
    equaln #(12) e2249(.a(buffered_input), .b(12'b100011001001), .eq(weq2249));
    equaln #(12) e2250(.a(buffered_input), .b(12'b100011001010), .eq(weq2250));
    equaln #(12) e2251(.a(buffered_input), .b(12'b100011001011), .eq(weq2251));
    equaln #(12) e2252(.a(buffered_input), .b(12'b100011001100), .eq(weq2252));
    equaln #(12) e2253(.a(buffered_input), .b(12'b100011001101), .eq(weq2253));
    equaln #(12) e2254(.a(buffered_input), .b(12'b100011001110), .eq(weq2254));
    equaln #(12) e2255(.a(buffered_input), .b(12'b100011001111), .eq(weq2255));
    equaln #(12) e2256(.a(buffered_input), .b(12'b100011010000), .eq(weq2256));
    equaln #(12) e2257(.a(buffered_input), .b(12'b100011010001), .eq(weq2257));
    equaln #(12) e2258(.a(buffered_input), .b(12'b100011010010), .eq(weq2258));
    equaln #(12) e2259(.a(buffered_input), .b(12'b100011010011), .eq(weq2259));
    equaln #(12) e2260(.a(buffered_input), .b(12'b100011010100), .eq(weq2260));
    equaln #(12) e2261(.a(buffered_input), .b(12'b100011010101), .eq(weq2261));
    equaln #(12) e2262(.a(buffered_input), .b(12'b100011010110), .eq(weq2262));
    equaln #(12) e2263(.a(buffered_input), .b(12'b100011010111), .eq(weq2263));
    equaln #(12) e2264(.a(buffered_input), .b(12'b100011011000), .eq(weq2264));
    equaln #(12) e2265(.a(buffered_input), .b(12'b100011011001), .eq(weq2265));
    equaln #(12) e2266(.a(buffered_input), .b(12'b100011011010), .eq(weq2266));
    equaln #(12) e2267(.a(buffered_input), .b(12'b100011011011), .eq(weq2267));
    equaln #(12) e2268(.a(buffered_input), .b(12'b100011011100), .eq(weq2268));
    equaln #(12) e2269(.a(buffered_input), .b(12'b100011011101), .eq(weq2269));
    equaln #(12) e2270(.a(buffered_input), .b(12'b100011011110), .eq(weq2270));
    equaln #(12) e2271(.a(buffered_input), .b(12'b100011011111), .eq(weq2271));
    equaln #(12) e2272(.a(buffered_input), .b(12'b100011100000), .eq(weq2272));
    equaln #(12) e2273(.a(buffered_input), .b(12'b100011100001), .eq(weq2273));
    equaln #(12) e2274(.a(buffered_input), .b(12'b100011100010), .eq(weq2274));
    equaln #(12) e2275(.a(buffered_input), .b(12'b100011100011), .eq(weq2275));
    equaln #(12) e2276(.a(buffered_input), .b(12'b100011100100), .eq(weq2276));
    equaln #(12) e2277(.a(buffered_input), .b(12'b100011100101), .eq(weq2277));
    equaln #(12) e2278(.a(buffered_input), .b(12'b100011100110), .eq(weq2278));
    equaln #(12) e2279(.a(buffered_input), .b(12'b100011100111), .eq(weq2279));
    equaln #(12) e2280(.a(buffered_input), .b(12'b100011101000), .eq(weq2280));
    equaln #(12) e2281(.a(buffered_input), .b(12'b100011101001), .eq(weq2281));
    equaln #(12) e2282(.a(buffered_input), .b(12'b100011101010), .eq(weq2282));
    equaln #(12) e2283(.a(buffered_input), .b(12'b100011101011), .eq(weq2283));
    equaln #(12) e2284(.a(buffered_input), .b(12'b100011101100), .eq(weq2284));
    equaln #(12) e2285(.a(buffered_input), .b(12'b100011101101), .eq(weq2285));
    equaln #(12) e2286(.a(buffered_input), .b(12'b100011101110), .eq(weq2286));
    equaln #(12) e2287(.a(buffered_input), .b(12'b100011101111), .eq(weq2287));
    equaln #(12) e2288(.a(buffered_input), .b(12'b100011110000), .eq(weq2288));
    equaln #(12) e2289(.a(buffered_input), .b(12'b100011110001), .eq(weq2289));
    equaln #(12) e2290(.a(buffered_input), .b(12'b100011110010), .eq(weq2290));
    equaln #(12) e2291(.a(buffered_input), .b(12'b100011110011), .eq(weq2291));
    equaln #(12) e2292(.a(buffered_input), .b(12'b100011110100), .eq(weq2292));
    equaln #(12) e2293(.a(buffered_input), .b(12'b100011110101), .eq(weq2293));
    equaln #(12) e2294(.a(buffered_input), .b(12'b100011110110), .eq(weq2294));
    equaln #(12) e2295(.a(buffered_input), .b(12'b100011110111), .eq(weq2295));
    equaln #(12) e2296(.a(buffered_input), .b(12'b100011111000), .eq(weq2296));
    equaln #(12) e2297(.a(buffered_input), .b(12'b100011111001), .eq(weq2297));
    equaln #(12) e2298(.a(buffered_input), .b(12'b100011111010), .eq(weq2298));
    equaln #(12) e2299(.a(buffered_input), .b(12'b100011111011), .eq(weq2299));
    equaln #(12) e2300(.a(buffered_input), .b(12'b100011111100), .eq(weq2300));
    equaln #(12) e2301(.a(buffered_input), .b(12'b100011111101), .eq(weq2301));
    equaln #(12) e2302(.a(buffered_input), .b(12'b100011111110), .eq(weq2302));
    equaln #(12) e2303(.a(buffered_input), .b(12'b100011111111), .eq(weq2303));
    equaln #(12) e2304(.a(buffered_input), .b(12'b100100000000), .eq(weq2304));
    equaln #(12) e2305(.a(buffered_input), .b(12'b100100000001), .eq(weq2305));
    equaln #(12) e2306(.a(buffered_input), .b(12'b100100000010), .eq(weq2306));
    equaln #(12) e2307(.a(buffered_input), .b(12'b100100000011), .eq(weq2307));
    equaln #(12) e2308(.a(buffered_input), .b(12'b100100000100), .eq(weq2308));
    equaln #(12) e2309(.a(buffered_input), .b(12'b100100000101), .eq(weq2309));
    equaln #(12) e2310(.a(buffered_input), .b(12'b100100000110), .eq(weq2310));
    equaln #(12) e2311(.a(buffered_input), .b(12'b100100000111), .eq(weq2311));
    equaln #(12) e2312(.a(buffered_input), .b(12'b100100001000), .eq(weq2312));
    equaln #(12) e2313(.a(buffered_input), .b(12'b100100001001), .eq(weq2313));
    equaln #(12) e2314(.a(buffered_input), .b(12'b100100001010), .eq(weq2314));
    equaln #(12) e2315(.a(buffered_input), .b(12'b100100001011), .eq(weq2315));
    equaln #(12) e2316(.a(buffered_input), .b(12'b100100001100), .eq(weq2316));
    equaln #(12) e2317(.a(buffered_input), .b(12'b100100001101), .eq(weq2317));
    equaln #(12) e2318(.a(buffered_input), .b(12'b100100001110), .eq(weq2318));
    equaln #(12) e2319(.a(buffered_input), .b(12'b100100001111), .eq(weq2319));
    equaln #(12) e2320(.a(buffered_input), .b(12'b100100010000), .eq(weq2320));
    equaln #(12) e2321(.a(buffered_input), .b(12'b100100010001), .eq(weq2321));
    equaln #(12) e2322(.a(buffered_input), .b(12'b100100010010), .eq(weq2322));
    equaln #(12) e2323(.a(buffered_input), .b(12'b100100010011), .eq(weq2323));
    equaln #(12) e2324(.a(buffered_input), .b(12'b100100010100), .eq(weq2324));
    equaln #(12) e2325(.a(buffered_input), .b(12'b100100010101), .eq(weq2325));
    equaln #(12) e2326(.a(buffered_input), .b(12'b100100010110), .eq(weq2326));
    equaln #(12) e2327(.a(buffered_input), .b(12'b100100010111), .eq(weq2327));
    equaln #(12) e2328(.a(buffered_input), .b(12'b100100011000), .eq(weq2328));
    equaln #(12) e2329(.a(buffered_input), .b(12'b100100011001), .eq(weq2329));
    equaln #(12) e2330(.a(buffered_input), .b(12'b100100011010), .eq(weq2330));
    equaln #(12) e2331(.a(buffered_input), .b(12'b100100011011), .eq(weq2331));
    equaln #(12) e2332(.a(buffered_input), .b(12'b100100011100), .eq(weq2332));
    equaln #(12) e2333(.a(buffered_input), .b(12'b100100011101), .eq(weq2333));
    equaln #(12) e2334(.a(buffered_input), .b(12'b100100011110), .eq(weq2334));
    equaln #(12) e2335(.a(buffered_input), .b(12'b100100011111), .eq(weq2335));
    equaln #(12) e2336(.a(buffered_input), .b(12'b100100100000), .eq(weq2336));
    equaln #(12) e2337(.a(buffered_input), .b(12'b100100100001), .eq(weq2337));
    equaln #(12) e2338(.a(buffered_input), .b(12'b100100100010), .eq(weq2338));
    equaln #(12) e2339(.a(buffered_input), .b(12'b100100100011), .eq(weq2339));
    equaln #(12) e2340(.a(buffered_input), .b(12'b100100100100), .eq(weq2340));
    equaln #(12) e2341(.a(buffered_input), .b(12'b100100100101), .eq(weq2341));
    equaln #(12) e2342(.a(buffered_input), .b(12'b100100100110), .eq(weq2342));
    equaln #(12) e2343(.a(buffered_input), .b(12'b100100100111), .eq(weq2343));
    equaln #(12) e2344(.a(buffered_input), .b(12'b100100101000), .eq(weq2344));
    equaln #(12) e2345(.a(buffered_input), .b(12'b100100101001), .eq(weq2345));
    equaln #(12) e2346(.a(buffered_input), .b(12'b100100101010), .eq(weq2346));
    equaln #(12) e2347(.a(buffered_input), .b(12'b100100101011), .eq(weq2347));
    equaln #(12) e2348(.a(buffered_input), .b(12'b100100101100), .eq(weq2348));
    equaln #(12) e2349(.a(buffered_input), .b(12'b100100101101), .eq(weq2349));
    equaln #(12) e2350(.a(buffered_input), .b(12'b100100101110), .eq(weq2350));
    equaln #(12) e2351(.a(buffered_input), .b(12'b100100101111), .eq(weq2351));
    equaln #(12) e2352(.a(buffered_input), .b(12'b100100110000), .eq(weq2352));
    equaln #(12) e2353(.a(buffered_input), .b(12'b100100110001), .eq(weq2353));
    equaln #(12) e2354(.a(buffered_input), .b(12'b100100110010), .eq(weq2354));
    equaln #(12) e2355(.a(buffered_input), .b(12'b100100110011), .eq(weq2355));
    equaln #(12) e2356(.a(buffered_input), .b(12'b100100110100), .eq(weq2356));
    equaln #(12) e2357(.a(buffered_input), .b(12'b100100110101), .eq(weq2357));
    equaln #(12) e2358(.a(buffered_input), .b(12'b100100110110), .eq(weq2358));
    equaln #(12) e2359(.a(buffered_input), .b(12'b100100110111), .eq(weq2359));
    equaln #(12) e2360(.a(buffered_input), .b(12'b100100111000), .eq(weq2360));
    equaln #(12) e2361(.a(buffered_input), .b(12'b100100111001), .eq(weq2361));
    equaln #(12) e2362(.a(buffered_input), .b(12'b100100111010), .eq(weq2362));
    equaln #(12) e2363(.a(buffered_input), .b(12'b100100111011), .eq(weq2363));
    equaln #(12) e2364(.a(buffered_input), .b(12'b100100111100), .eq(weq2364));
    equaln #(12) e2365(.a(buffered_input), .b(12'b100100111101), .eq(weq2365));
    equaln #(12) e2366(.a(buffered_input), .b(12'b100100111110), .eq(weq2366));
    equaln #(12) e2367(.a(buffered_input), .b(12'b100100111111), .eq(weq2367));
    equaln #(12) e2368(.a(buffered_input), .b(12'b100101000000), .eq(weq2368));
    equaln #(12) e2369(.a(buffered_input), .b(12'b100101000001), .eq(weq2369));
    equaln #(12) e2370(.a(buffered_input), .b(12'b100101000010), .eq(weq2370));
    equaln #(12) e2371(.a(buffered_input), .b(12'b100101000011), .eq(weq2371));
    equaln #(12) e2372(.a(buffered_input), .b(12'b100101000100), .eq(weq2372));
    equaln #(12) e2373(.a(buffered_input), .b(12'b100101000101), .eq(weq2373));
    equaln #(12) e2374(.a(buffered_input), .b(12'b100101000110), .eq(weq2374));
    equaln #(12) e2375(.a(buffered_input), .b(12'b100101000111), .eq(weq2375));
    equaln #(12) e2376(.a(buffered_input), .b(12'b100101001000), .eq(weq2376));
    equaln #(12) e2377(.a(buffered_input), .b(12'b100101001001), .eq(weq2377));
    equaln #(12) e2378(.a(buffered_input), .b(12'b100101001010), .eq(weq2378));
    equaln #(12) e2379(.a(buffered_input), .b(12'b100101001011), .eq(weq2379));
    equaln #(12) e2380(.a(buffered_input), .b(12'b100101001100), .eq(weq2380));
    equaln #(12) e2381(.a(buffered_input), .b(12'b100101001101), .eq(weq2381));
    equaln #(12) e2382(.a(buffered_input), .b(12'b100101001110), .eq(weq2382));
    equaln #(12) e2383(.a(buffered_input), .b(12'b100101001111), .eq(weq2383));
    equaln #(12) e2384(.a(buffered_input), .b(12'b100101010000), .eq(weq2384));
    equaln #(12) e2385(.a(buffered_input), .b(12'b100101010001), .eq(weq2385));
    equaln #(12) e2386(.a(buffered_input), .b(12'b100101010010), .eq(weq2386));
    equaln #(12) e2387(.a(buffered_input), .b(12'b100101010011), .eq(weq2387));
    equaln #(12) e2388(.a(buffered_input), .b(12'b100101010100), .eq(weq2388));
    equaln #(12) e2389(.a(buffered_input), .b(12'b100101010101), .eq(weq2389));
    equaln #(12) e2390(.a(buffered_input), .b(12'b100101010110), .eq(weq2390));
    equaln #(12) e2391(.a(buffered_input), .b(12'b100101010111), .eq(weq2391));
    equaln #(12) e2392(.a(buffered_input), .b(12'b100101011000), .eq(weq2392));
    equaln #(12) e2393(.a(buffered_input), .b(12'b100101011001), .eq(weq2393));
    equaln #(12) e2394(.a(buffered_input), .b(12'b100101011010), .eq(weq2394));
    equaln #(12) e2395(.a(buffered_input), .b(12'b100101011011), .eq(weq2395));
    equaln #(12) e2396(.a(buffered_input), .b(12'b100101011100), .eq(weq2396));
    equaln #(12) e2397(.a(buffered_input), .b(12'b100101011101), .eq(weq2397));
    equaln #(12) e2398(.a(buffered_input), .b(12'b100101011110), .eq(weq2398));
    equaln #(12) e2399(.a(buffered_input), .b(12'b100101011111), .eq(weq2399));
    equaln #(12) e2400(.a(buffered_input), .b(12'b100101100000), .eq(weq2400));
    equaln #(12) e2401(.a(buffered_input), .b(12'b100101100001), .eq(weq2401));
    equaln #(12) e2402(.a(buffered_input), .b(12'b100101100010), .eq(weq2402));
    equaln #(12) e2403(.a(buffered_input), .b(12'b100101100011), .eq(weq2403));
    equaln #(12) e2404(.a(buffered_input), .b(12'b100101100100), .eq(weq2404));
    equaln #(12) e2405(.a(buffered_input), .b(12'b100101100101), .eq(weq2405));
    equaln #(12) e2406(.a(buffered_input), .b(12'b100101100110), .eq(weq2406));
    equaln #(12) e2407(.a(buffered_input), .b(12'b100101100111), .eq(weq2407));
    equaln #(12) e2408(.a(buffered_input), .b(12'b100101101000), .eq(weq2408));
    equaln #(12) e2409(.a(buffered_input), .b(12'b100101101001), .eq(weq2409));
    equaln #(12) e2410(.a(buffered_input), .b(12'b100101101010), .eq(weq2410));
    equaln #(12) e2411(.a(buffered_input), .b(12'b100101101011), .eq(weq2411));
    equaln #(12) e2412(.a(buffered_input), .b(12'b100101101100), .eq(weq2412));
    equaln #(12) e2413(.a(buffered_input), .b(12'b100101101101), .eq(weq2413));
    equaln #(12) e2414(.a(buffered_input), .b(12'b100101101110), .eq(weq2414));
    equaln #(12) e2415(.a(buffered_input), .b(12'b100101101111), .eq(weq2415));
    equaln #(12) e2416(.a(buffered_input), .b(12'b100101110000), .eq(weq2416));
    equaln #(12) e2417(.a(buffered_input), .b(12'b100101110001), .eq(weq2417));
    equaln #(12) e2418(.a(buffered_input), .b(12'b100101110010), .eq(weq2418));
    equaln #(12) e2419(.a(buffered_input), .b(12'b100101110011), .eq(weq2419));
    equaln #(12) e2420(.a(buffered_input), .b(12'b100101110100), .eq(weq2420));
    equaln #(12) e2421(.a(buffered_input), .b(12'b100101110101), .eq(weq2421));
    equaln #(12) e2422(.a(buffered_input), .b(12'b100101110110), .eq(weq2422));
    equaln #(12) e2423(.a(buffered_input), .b(12'b100101110111), .eq(weq2423));
    equaln #(12) e2424(.a(buffered_input), .b(12'b100101111000), .eq(weq2424));
    equaln #(12) e2425(.a(buffered_input), .b(12'b100101111001), .eq(weq2425));
    equaln #(12) e2426(.a(buffered_input), .b(12'b100101111010), .eq(weq2426));
    equaln #(12) e2427(.a(buffered_input), .b(12'b100101111011), .eq(weq2427));
    equaln #(12) e2428(.a(buffered_input), .b(12'b100101111100), .eq(weq2428));
    equaln #(12) e2429(.a(buffered_input), .b(12'b100101111101), .eq(weq2429));
    equaln #(12) e2430(.a(buffered_input), .b(12'b100101111110), .eq(weq2430));
    equaln #(12) e2431(.a(buffered_input), .b(12'b100101111111), .eq(weq2431));
    equaln #(12) e2432(.a(buffered_input), .b(12'b100110000000), .eq(weq2432));
    equaln #(12) e2433(.a(buffered_input), .b(12'b100110000001), .eq(weq2433));
    equaln #(12) e2434(.a(buffered_input), .b(12'b100110000010), .eq(weq2434));
    equaln #(12) e2435(.a(buffered_input), .b(12'b100110000011), .eq(weq2435));
    equaln #(12) e2436(.a(buffered_input), .b(12'b100110000100), .eq(weq2436));
    equaln #(12) e2437(.a(buffered_input), .b(12'b100110000101), .eq(weq2437));
    equaln #(12) e2438(.a(buffered_input), .b(12'b100110000110), .eq(weq2438));
    equaln #(12) e2439(.a(buffered_input), .b(12'b100110000111), .eq(weq2439));
    equaln #(12) e2440(.a(buffered_input), .b(12'b100110001000), .eq(weq2440));
    equaln #(12) e2441(.a(buffered_input), .b(12'b100110001001), .eq(weq2441));
    equaln #(12) e2442(.a(buffered_input), .b(12'b100110001010), .eq(weq2442));
    equaln #(12) e2443(.a(buffered_input), .b(12'b100110001011), .eq(weq2443));
    equaln #(12) e2444(.a(buffered_input), .b(12'b100110001100), .eq(weq2444));
    equaln #(12) e2445(.a(buffered_input), .b(12'b100110001101), .eq(weq2445));
    equaln #(12) e2446(.a(buffered_input), .b(12'b100110001110), .eq(weq2446));
    equaln #(12) e2447(.a(buffered_input), .b(12'b100110001111), .eq(weq2447));
    equaln #(12) e2448(.a(buffered_input), .b(12'b100110010000), .eq(weq2448));
    equaln #(12) e2449(.a(buffered_input), .b(12'b100110010001), .eq(weq2449));
    equaln #(12) e2450(.a(buffered_input), .b(12'b100110010010), .eq(weq2450));
    equaln #(12) e2451(.a(buffered_input), .b(12'b100110010011), .eq(weq2451));
    equaln #(12) e2452(.a(buffered_input), .b(12'b100110010100), .eq(weq2452));
    equaln #(12) e2453(.a(buffered_input), .b(12'b100110010101), .eq(weq2453));
    equaln #(12) e2454(.a(buffered_input), .b(12'b100110010110), .eq(weq2454));
    equaln #(12) e2455(.a(buffered_input), .b(12'b100110010111), .eq(weq2455));
    equaln #(12) e2456(.a(buffered_input), .b(12'b100110011000), .eq(weq2456));
    equaln #(12) e2457(.a(buffered_input), .b(12'b100110011001), .eq(weq2457));
    equaln #(12) e2458(.a(buffered_input), .b(12'b100110011010), .eq(weq2458));
    equaln #(12) e2459(.a(buffered_input), .b(12'b100110011011), .eq(weq2459));
    equaln #(12) e2460(.a(buffered_input), .b(12'b100110011100), .eq(weq2460));
    equaln #(12) e2461(.a(buffered_input), .b(12'b100110011101), .eq(weq2461));
    equaln #(12) e2462(.a(buffered_input), .b(12'b100110011110), .eq(weq2462));
    equaln #(12) e2463(.a(buffered_input), .b(12'b100110011111), .eq(weq2463));
    equaln #(12) e2464(.a(buffered_input), .b(12'b100110100000), .eq(weq2464));
    equaln #(12) e2465(.a(buffered_input), .b(12'b100110100001), .eq(weq2465));
    equaln #(12) e2466(.a(buffered_input), .b(12'b100110100010), .eq(weq2466));
    equaln #(12) e2467(.a(buffered_input), .b(12'b100110100011), .eq(weq2467));
    equaln #(12) e2468(.a(buffered_input), .b(12'b100110100100), .eq(weq2468));
    equaln #(12) e2469(.a(buffered_input), .b(12'b100110100101), .eq(weq2469));
    equaln #(12) e2470(.a(buffered_input), .b(12'b100110100110), .eq(weq2470));
    equaln #(12) e2471(.a(buffered_input), .b(12'b100110100111), .eq(weq2471));
    equaln #(12) e2472(.a(buffered_input), .b(12'b100110101000), .eq(weq2472));
    equaln #(12) e2473(.a(buffered_input), .b(12'b100110101001), .eq(weq2473));
    equaln #(12) e2474(.a(buffered_input), .b(12'b100110101010), .eq(weq2474));
    equaln #(12) e2475(.a(buffered_input), .b(12'b100110101011), .eq(weq2475));
    equaln #(12) e2476(.a(buffered_input), .b(12'b100110101100), .eq(weq2476));
    equaln #(12) e2477(.a(buffered_input), .b(12'b100110101101), .eq(weq2477));
    equaln #(12) e2478(.a(buffered_input), .b(12'b100110101110), .eq(weq2478));
    equaln #(12) e2479(.a(buffered_input), .b(12'b100110101111), .eq(weq2479));
    equaln #(12) e2480(.a(buffered_input), .b(12'b100110110000), .eq(weq2480));
    equaln #(12) e2481(.a(buffered_input), .b(12'b100110110001), .eq(weq2481));
    equaln #(12) e2482(.a(buffered_input), .b(12'b100110110010), .eq(weq2482));
    equaln #(12) e2483(.a(buffered_input), .b(12'b100110110011), .eq(weq2483));
    equaln #(12) e2484(.a(buffered_input), .b(12'b100110110100), .eq(weq2484));
    equaln #(12) e2485(.a(buffered_input), .b(12'b100110110101), .eq(weq2485));
    equaln #(12) e2486(.a(buffered_input), .b(12'b100110110110), .eq(weq2486));
    equaln #(12) e2487(.a(buffered_input), .b(12'b100110110111), .eq(weq2487));
    equaln #(12) e2488(.a(buffered_input), .b(12'b100110111000), .eq(weq2488));
    equaln #(12) e2489(.a(buffered_input), .b(12'b100110111001), .eq(weq2489));
    equaln #(12) e2490(.a(buffered_input), .b(12'b100110111010), .eq(weq2490));
    equaln #(12) e2491(.a(buffered_input), .b(12'b100110111011), .eq(weq2491));
    equaln #(12) e2492(.a(buffered_input), .b(12'b100110111100), .eq(weq2492));
    equaln #(12) e2493(.a(buffered_input), .b(12'b100110111101), .eq(weq2493));
    equaln #(12) e2494(.a(buffered_input), .b(12'b100110111110), .eq(weq2494));
    equaln #(12) e2495(.a(buffered_input), .b(12'b100110111111), .eq(weq2495));
    equaln #(12) e2496(.a(buffered_input), .b(12'b100111000000), .eq(weq2496));
    equaln #(12) e2497(.a(buffered_input), .b(12'b100111000001), .eq(weq2497));
    equaln #(12) e2498(.a(buffered_input), .b(12'b100111000010), .eq(weq2498));
    equaln #(12) e2499(.a(buffered_input), .b(12'b100111000011), .eq(weq2499));
    equaln #(12) e2500(.a(buffered_input), .b(12'b100111000100), .eq(weq2500));
    equaln #(12) e2501(.a(buffered_input), .b(12'b100111000101), .eq(weq2501));
    equaln #(12) e2502(.a(buffered_input), .b(12'b100111000110), .eq(weq2502));
    equaln #(12) e2503(.a(buffered_input), .b(12'b100111000111), .eq(weq2503));
    equaln #(12) e2504(.a(buffered_input), .b(12'b100111001000), .eq(weq2504));
    equaln #(12) e2505(.a(buffered_input), .b(12'b100111001001), .eq(weq2505));
    equaln #(12) e2506(.a(buffered_input), .b(12'b100111001010), .eq(weq2506));
    equaln #(12) e2507(.a(buffered_input), .b(12'b100111001011), .eq(weq2507));
    equaln #(12) e2508(.a(buffered_input), .b(12'b100111001100), .eq(weq2508));
    equaln #(12) e2509(.a(buffered_input), .b(12'b100111001101), .eq(weq2509));
    equaln #(12) e2510(.a(buffered_input), .b(12'b100111001110), .eq(weq2510));
    equaln #(12) e2511(.a(buffered_input), .b(12'b100111001111), .eq(weq2511));
    equaln #(12) e2512(.a(buffered_input), .b(12'b100111010000), .eq(weq2512));
    equaln #(12) e2513(.a(buffered_input), .b(12'b100111010001), .eq(weq2513));
    equaln #(12) e2514(.a(buffered_input), .b(12'b100111010010), .eq(weq2514));
    equaln #(12) e2515(.a(buffered_input), .b(12'b100111010011), .eq(weq2515));
    equaln #(12) e2516(.a(buffered_input), .b(12'b100111010100), .eq(weq2516));
    equaln #(12) e2517(.a(buffered_input), .b(12'b100111010101), .eq(weq2517));
    equaln #(12) e2518(.a(buffered_input), .b(12'b100111010110), .eq(weq2518));
    equaln #(12) e2519(.a(buffered_input), .b(12'b100111010111), .eq(weq2519));
    equaln #(12) e2520(.a(buffered_input), .b(12'b100111011000), .eq(weq2520));
    equaln #(12) e2521(.a(buffered_input), .b(12'b100111011001), .eq(weq2521));
    equaln #(12) e2522(.a(buffered_input), .b(12'b100111011010), .eq(weq2522));
    equaln #(12) e2523(.a(buffered_input), .b(12'b100111011011), .eq(weq2523));
    equaln #(12) e2524(.a(buffered_input), .b(12'b100111011100), .eq(weq2524));
    equaln #(12) e2525(.a(buffered_input), .b(12'b100111011101), .eq(weq2525));
    equaln #(12) e2526(.a(buffered_input), .b(12'b100111011110), .eq(weq2526));
    equaln #(12) e2527(.a(buffered_input), .b(12'b100111011111), .eq(weq2527));
    equaln #(12) e2528(.a(buffered_input), .b(12'b100111100000), .eq(weq2528));
    equaln #(12) e2529(.a(buffered_input), .b(12'b100111100001), .eq(weq2529));
    equaln #(12) e2530(.a(buffered_input), .b(12'b100111100010), .eq(weq2530));
    equaln #(12) e2531(.a(buffered_input), .b(12'b100111100011), .eq(weq2531));
    equaln #(12) e2532(.a(buffered_input), .b(12'b100111100100), .eq(weq2532));
    equaln #(12) e2533(.a(buffered_input), .b(12'b100111100101), .eq(weq2533));
    equaln #(12) e2534(.a(buffered_input), .b(12'b100111100110), .eq(weq2534));
    equaln #(12) e2535(.a(buffered_input), .b(12'b100111100111), .eq(weq2535));
    equaln #(12) e2536(.a(buffered_input), .b(12'b100111101000), .eq(weq2536));
    equaln #(12) e2537(.a(buffered_input), .b(12'b100111101001), .eq(weq2537));
    equaln #(12) e2538(.a(buffered_input), .b(12'b100111101010), .eq(weq2538));
    equaln #(12) e2539(.a(buffered_input), .b(12'b100111101011), .eq(weq2539));
    equaln #(12) e2540(.a(buffered_input), .b(12'b100111101100), .eq(weq2540));
    equaln #(12) e2541(.a(buffered_input), .b(12'b100111101101), .eq(weq2541));
    equaln #(12) e2542(.a(buffered_input), .b(12'b100111101110), .eq(weq2542));
    equaln #(12) e2543(.a(buffered_input), .b(12'b100111101111), .eq(weq2543));
    equaln #(12) e2544(.a(buffered_input), .b(12'b100111110000), .eq(weq2544));
    equaln #(12) e2545(.a(buffered_input), .b(12'b100111110001), .eq(weq2545));
    equaln #(12) e2546(.a(buffered_input), .b(12'b100111110010), .eq(weq2546));
    equaln #(12) e2547(.a(buffered_input), .b(12'b100111110011), .eq(weq2547));
    equaln #(12) e2548(.a(buffered_input), .b(12'b100111110100), .eq(weq2548));
    equaln #(12) e2549(.a(buffered_input), .b(12'b100111110101), .eq(weq2549));
    equaln #(12) e2550(.a(buffered_input), .b(12'b100111110110), .eq(weq2550));
    equaln #(12) e2551(.a(buffered_input), .b(12'b100111110111), .eq(weq2551));
    equaln #(12) e2552(.a(buffered_input), .b(12'b100111111000), .eq(weq2552));
    equaln #(12) e2553(.a(buffered_input), .b(12'b100111111001), .eq(weq2553));
    equaln #(12) e2554(.a(buffered_input), .b(12'b100111111010), .eq(weq2554));
    equaln #(12) e2555(.a(buffered_input), .b(12'b100111111011), .eq(weq2555));
    equaln #(12) e2556(.a(buffered_input), .b(12'b100111111100), .eq(weq2556));
    equaln #(12) e2557(.a(buffered_input), .b(12'b100111111101), .eq(weq2557));
    equaln #(12) e2558(.a(buffered_input), .b(12'b100111111110), .eq(weq2558));
    equaln #(12) e2559(.a(buffered_input), .b(12'b100111111111), .eq(weq2559));
    equaln #(12) e2560(.a(buffered_input), .b(12'b101000000000), .eq(weq2560));
    equaln #(12) e2561(.a(buffered_input), .b(12'b101000000001), .eq(weq2561));
    equaln #(12) e2562(.a(buffered_input), .b(12'b101000000010), .eq(weq2562));
    equaln #(12) e2563(.a(buffered_input), .b(12'b101000000011), .eq(weq2563));
    equaln #(12) e2564(.a(buffered_input), .b(12'b101000000100), .eq(weq2564));
    equaln #(12) e2565(.a(buffered_input), .b(12'b101000000101), .eq(weq2565));
    equaln #(12) e2566(.a(buffered_input), .b(12'b101000000110), .eq(weq2566));
    equaln #(12) e2567(.a(buffered_input), .b(12'b101000000111), .eq(weq2567));
    equaln #(12) e2568(.a(buffered_input), .b(12'b101000001000), .eq(weq2568));
    equaln #(12) e2569(.a(buffered_input), .b(12'b101000001001), .eq(weq2569));
    equaln #(12) e2570(.a(buffered_input), .b(12'b101000001010), .eq(weq2570));
    equaln #(12) e2571(.a(buffered_input), .b(12'b101000001011), .eq(weq2571));
    equaln #(12) e2572(.a(buffered_input), .b(12'b101000001100), .eq(weq2572));
    equaln #(12) e2573(.a(buffered_input), .b(12'b101000001101), .eq(weq2573));
    equaln #(12) e2574(.a(buffered_input), .b(12'b101000001110), .eq(weq2574));
    equaln #(12) e2575(.a(buffered_input), .b(12'b101000001111), .eq(weq2575));
    equaln #(12) e2576(.a(buffered_input), .b(12'b101000010000), .eq(weq2576));
    equaln #(12) e2577(.a(buffered_input), .b(12'b101000010001), .eq(weq2577));
    equaln #(12) e2578(.a(buffered_input), .b(12'b101000010010), .eq(weq2578));
    equaln #(12) e2579(.a(buffered_input), .b(12'b101000010011), .eq(weq2579));
    equaln #(12) e2580(.a(buffered_input), .b(12'b101000010100), .eq(weq2580));
    equaln #(12) e2581(.a(buffered_input), .b(12'b101000010101), .eq(weq2581));
    equaln #(12) e2582(.a(buffered_input), .b(12'b101000010110), .eq(weq2582));
    equaln #(12) e2583(.a(buffered_input), .b(12'b101000010111), .eq(weq2583));
    equaln #(12) e2584(.a(buffered_input), .b(12'b101000011000), .eq(weq2584));
    equaln #(12) e2585(.a(buffered_input), .b(12'b101000011001), .eq(weq2585));
    equaln #(12) e2586(.a(buffered_input), .b(12'b101000011010), .eq(weq2586));
    equaln #(12) e2587(.a(buffered_input), .b(12'b101000011011), .eq(weq2587));
    equaln #(12) e2588(.a(buffered_input), .b(12'b101000011100), .eq(weq2588));
    equaln #(12) e2589(.a(buffered_input), .b(12'b101000011101), .eq(weq2589));
    equaln #(12) e2590(.a(buffered_input), .b(12'b101000011110), .eq(weq2590));
    equaln #(12) e2591(.a(buffered_input), .b(12'b101000011111), .eq(weq2591));
    equaln #(12) e2592(.a(buffered_input), .b(12'b101000100000), .eq(weq2592));
    equaln #(12) e2593(.a(buffered_input), .b(12'b101000100001), .eq(weq2593));
    equaln #(12) e2594(.a(buffered_input), .b(12'b101000100010), .eq(weq2594));
    equaln #(12) e2595(.a(buffered_input), .b(12'b101000100011), .eq(weq2595));
    equaln #(12) e2596(.a(buffered_input), .b(12'b101000100100), .eq(weq2596));
    equaln #(12) e2597(.a(buffered_input), .b(12'b101000100101), .eq(weq2597));
    equaln #(12) e2598(.a(buffered_input), .b(12'b101000100110), .eq(weq2598));
    equaln #(12) e2599(.a(buffered_input), .b(12'b101000100111), .eq(weq2599));
    equaln #(12) e2600(.a(buffered_input), .b(12'b101000101000), .eq(weq2600));
    equaln #(12) e2601(.a(buffered_input), .b(12'b101000101001), .eq(weq2601));
    equaln #(12) e2602(.a(buffered_input), .b(12'b101000101010), .eq(weq2602));
    equaln #(12) e2603(.a(buffered_input), .b(12'b101000101011), .eq(weq2603));
    equaln #(12) e2604(.a(buffered_input), .b(12'b101000101100), .eq(weq2604));
    equaln #(12) e2605(.a(buffered_input), .b(12'b101000101101), .eq(weq2605));
    equaln #(12) e2606(.a(buffered_input), .b(12'b101000101110), .eq(weq2606));
    equaln #(12) e2607(.a(buffered_input), .b(12'b101000101111), .eq(weq2607));
    equaln #(12) e2608(.a(buffered_input), .b(12'b101000110000), .eq(weq2608));
    equaln #(12) e2609(.a(buffered_input), .b(12'b101000110001), .eq(weq2609));
    equaln #(12) e2610(.a(buffered_input), .b(12'b101000110010), .eq(weq2610));
    equaln #(12) e2611(.a(buffered_input), .b(12'b101000110011), .eq(weq2611));
    equaln #(12) e2612(.a(buffered_input), .b(12'b101000110100), .eq(weq2612));
    equaln #(12) e2613(.a(buffered_input), .b(12'b101000110101), .eq(weq2613));
    equaln #(12) e2614(.a(buffered_input), .b(12'b101000110110), .eq(weq2614));
    equaln #(12) e2615(.a(buffered_input), .b(12'b101000110111), .eq(weq2615));
    equaln #(12) e2616(.a(buffered_input), .b(12'b101000111000), .eq(weq2616));
    equaln #(12) e2617(.a(buffered_input), .b(12'b101000111001), .eq(weq2617));
    equaln #(12) e2618(.a(buffered_input), .b(12'b101000111010), .eq(weq2618));
    equaln #(12) e2619(.a(buffered_input), .b(12'b101000111011), .eq(weq2619));
    equaln #(12) e2620(.a(buffered_input), .b(12'b101000111100), .eq(weq2620));
    equaln #(12) e2621(.a(buffered_input), .b(12'b101000111101), .eq(weq2621));
    equaln #(12) e2622(.a(buffered_input), .b(12'b101000111110), .eq(weq2622));
    equaln #(12) e2623(.a(buffered_input), .b(12'b101000111111), .eq(weq2623));
    equaln #(12) e2624(.a(buffered_input), .b(12'b101001000000), .eq(weq2624));
    equaln #(12) e2625(.a(buffered_input), .b(12'b101001000001), .eq(weq2625));
    equaln #(12) e2626(.a(buffered_input), .b(12'b101001000010), .eq(weq2626));
    equaln #(12) e2627(.a(buffered_input), .b(12'b101001000011), .eq(weq2627));
    equaln #(12) e2628(.a(buffered_input), .b(12'b101001000100), .eq(weq2628));
    equaln #(12) e2629(.a(buffered_input), .b(12'b101001000101), .eq(weq2629));
    equaln #(12) e2630(.a(buffered_input), .b(12'b101001000110), .eq(weq2630));
    equaln #(12) e2631(.a(buffered_input), .b(12'b101001000111), .eq(weq2631));
    equaln #(12) e2632(.a(buffered_input), .b(12'b101001001000), .eq(weq2632));
    equaln #(12) e2633(.a(buffered_input), .b(12'b101001001001), .eq(weq2633));
    equaln #(12) e2634(.a(buffered_input), .b(12'b101001001010), .eq(weq2634));
    equaln #(12) e2635(.a(buffered_input), .b(12'b101001001011), .eq(weq2635));
    equaln #(12) e2636(.a(buffered_input), .b(12'b101001001100), .eq(weq2636));
    equaln #(12) e2637(.a(buffered_input), .b(12'b101001001101), .eq(weq2637));
    equaln #(12) e2638(.a(buffered_input), .b(12'b101001001110), .eq(weq2638));
    equaln #(12) e2639(.a(buffered_input), .b(12'b101001001111), .eq(weq2639));
    equaln #(12) e2640(.a(buffered_input), .b(12'b101001010000), .eq(weq2640));
    equaln #(12) e2641(.a(buffered_input), .b(12'b101001010001), .eq(weq2641));
    equaln #(12) e2642(.a(buffered_input), .b(12'b101001010010), .eq(weq2642));
    equaln #(12) e2643(.a(buffered_input), .b(12'b101001010011), .eq(weq2643));
    equaln #(12) e2644(.a(buffered_input), .b(12'b101001010100), .eq(weq2644));
    equaln #(12) e2645(.a(buffered_input), .b(12'b101001010101), .eq(weq2645));
    equaln #(12) e2646(.a(buffered_input), .b(12'b101001010110), .eq(weq2646));
    equaln #(12) e2647(.a(buffered_input), .b(12'b101001010111), .eq(weq2647));
    equaln #(12) e2648(.a(buffered_input), .b(12'b101001011000), .eq(weq2648));
    equaln #(12) e2649(.a(buffered_input), .b(12'b101001011001), .eq(weq2649));
    equaln #(12) e2650(.a(buffered_input), .b(12'b101001011010), .eq(weq2650));
    equaln #(12) e2651(.a(buffered_input), .b(12'b101001011011), .eq(weq2651));
    equaln #(12) e2652(.a(buffered_input), .b(12'b101001011100), .eq(weq2652));
    equaln #(12) e2653(.a(buffered_input), .b(12'b101001011101), .eq(weq2653));
    equaln #(12) e2654(.a(buffered_input), .b(12'b101001011110), .eq(weq2654));
    equaln #(12) e2655(.a(buffered_input), .b(12'b101001011111), .eq(weq2655));
    equaln #(12) e2656(.a(buffered_input), .b(12'b101001100000), .eq(weq2656));
    equaln #(12) e2657(.a(buffered_input), .b(12'b101001100001), .eq(weq2657));
    equaln #(12) e2658(.a(buffered_input), .b(12'b101001100010), .eq(weq2658));
    equaln #(12) e2659(.a(buffered_input), .b(12'b101001100011), .eq(weq2659));
    equaln #(12) e2660(.a(buffered_input), .b(12'b101001100100), .eq(weq2660));
    equaln #(12) e2661(.a(buffered_input), .b(12'b101001100101), .eq(weq2661));
    equaln #(12) e2662(.a(buffered_input), .b(12'b101001100110), .eq(weq2662));
    equaln #(12) e2663(.a(buffered_input), .b(12'b101001100111), .eq(weq2663));
    equaln #(12) e2664(.a(buffered_input), .b(12'b101001101000), .eq(weq2664));
    equaln #(12) e2665(.a(buffered_input), .b(12'b101001101001), .eq(weq2665));
    equaln #(12) e2666(.a(buffered_input), .b(12'b101001101010), .eq(weq2666));
    equaln #(12) e2667(.a(buffered_input), .b(12'b101001101011), .eq(weq2667));
    equaln #(12) e2668(.a(buffered_input), .b(12'b101001101100), .eq(weq2668));
    equaln #(12) e2669(.a(buffered_input), .b(12'b101001101101), .eq(weq2669));
    equaln #(12) e2670(.a(buffered_input), .b(12'b101001101110), .eq(weq2670));
    equaln #(12) e2671(.a(buffered_input), .b(12'b101001101111), .eq(weq2671));
    equaln #(12) e2672(.a(buffered_input), .b(12'b101001110000), .eq(weq2672));
    equaln #(12) e2673(.a(buffered_input), .b(12'b101001110001), .eq(weq2673));
    equaln #(12) e2674(.a(buffered_input), .b(12'b101001110010), .eq(weq2674));
    equaln #(12) e2675(.a(buffered_input), .b(12'b101001110011), .eq(weq2675));
    equaln #(12) e2676(.a(buffered_input), .b(12'b101001110100), .eq(weq2676));
    equaln #(12) e2677(.a(buffered_input), .b(12'b101001110101), .eq(weq2677));
    equaln #(12) e2678(.a(buffered_input), .b(12'b101001110110), .eq(weq2678));
    equaln #(12) e2679(.a(buffered_input), .b(12'b101001110111), .eq(weq2679));
    equaln #(12) e2680(.a(buffered_input), .b(12'b101001111000), .eq(weq2680));
    equaln #(12) e2681(.a(buffered_input), .b(12'b101001111001), .eq(weq2681));
    equaln #(12) e2682(.a(buffered_input), .b(12'b101001111010), .eq(weq2682));
    equaln #(12) e2683(.a(buffered_input), .b(12'b101001111011), .eq(weq2683));
    equaln #(12) e2684(.a(buffered_input), .b(12'b101001111100), .eq(weq2684));
    equaln #(12) e2685(.a(buffered_input), .b(12'b101001111101), .eq(weq2685));
    equaln #(12) e2686(.a(buffered_input), .b(12'b101001111110), .eq(weq2686));
    equaln #(12) e2687(.a(buffered_input), .b(12'b101001111111), .eq(weq2687));
    equaln #(12) e2688(.a(buffered_input), .b(12'b101010000000), .eq(weq2688));
    equaln #(12) e2689(.a(buffered_input), .b(12'b101010000001), .eq(weq2689));
    equaln #(12) e2690(.a(buffered_input), .b(12'b101010000010), .eq(weq2690));
    equaln #(12) e2691(.a(buffered_input), .b(12'b101010000011), .eq(weq2691));
    equaln #(12) e2692(.a(buffered_input), .b(12'b101010000100), .eq(weq2692));
    equaln #(12) e2693(.a(buffered_input), .b(12'b101010000101), .eq(weq2693));
    equaln #(12) e2694(.a(buffered_input), .b(12'b101010000110), .eq(weq2694));
    equaln #(12) e2695(.a(buffered_input), .b(12'b101010000111), .eq(weq2695));
    equaln #(12) e2696(.a(buffered_input), .b(12'b101010001000), .eq(weq2696));
    equaln #(12) e2697(.a(buffered_input), .b(12'b101010001001), .eq(weq2697));
    equaln #(12) e2698(.a(buffered_input), .b(12'b101010001010), .eq(weq2698));
    equaln #(12) e2699(.a(buffered_input), .b(12'b101010001011), .eq(weq2699));
    equaln #(12) e2700(.a(buffered_input), .b(12'b101010001100), .eq(weq2700));
    equaln #(12) e2701(.a(buffered_input), .b(12'b101010001101), .eq(weq2701));
    equaln #(12) e2702(.a(buffered_input), .b(12'b101010001110), .eq(weq2702));
    equaln #(12) e2703(.a(buffered_input), .b(12'b101010001111), .eq(weq2703));
    equaln #(12) e2704(.a(buffered_input), .b(12'b101010010000), .eq(weq2704));
    equaln #(12) e2705(.a(buffered_input), .b(12'b101010010001), .eq(weq2705));
    equaln #(12) e2706(.a(buffered_input), .b(12'b101010010010), .eq(weq2706));
    equaln #(12) e2707(.a(buffered_input), .b(12'b101010010011), .eq(weq2707));
    equaln #(12) e2708(.a(buffered_input), .b(12'b101010010100), .eq(weq2708));
    equaln #(12) e2709(.a(buffered_input), .b(12'b101010010101), .eq(weq2709));
    equaln #(12) e2710(.a(buffered_input), .b(12'b101010010110), .eq(weq2710));
    equaln #(12) e2711(.a(buffered_input), .b(12'b101010010111), .eq(weq2711));
    equaln #(12) e2712(.a(buffered_input), .b(12'b101010011000), .eq(weq2712));
    equaln #(12) e2713(.a(buffered_input), .b(12'b101010011001), .eq(weq2713));
    equaln #(12) e2714(.a(buffered_input), .b(12'b101010011010), .eq(weq2714));
    equaln #(12) e2715(.a(buffered_input), .b(12'b101010011011), .eq(weq2715));
    equaln #(12) e2716(.a(buffered_input), .b(12'b101010011100), .eq(weq2716));
    equaln #(12) e2717(.a(buffered_input), .b(12'b101010011101), .eq(weq2717));
    equaln #(12) e2718(.a(buffered_input), .b(12'b101010011110), .eq(weq2718));
    equaln #(12) e2719(.a(buffered_input), .b(12'b101010011111), .eq(weq2719));
    equaln #(12) e2720(.a(buffered_input), .b(12'b101010100000), .eq(weq2720));
    equaln #(12) e2721(.a(buffered_input), .b(12'b101010100001), .eq(weq2721));
    equaln #(12) e2722(.a(buffered_input), .b(12'b101010100010), .eq(weq2722));
    equaln #(12) e2723(.a(buffered_input), .b(12'b101010100011), .eq(weq2723));
    equaln #(12) e2724(.a(buffered_input), .b(12'b101010100100), .eq(weq2724));
    equaln #(12) e2725(.a(buffered_input), .b(12'b101010100101), .eq(weq2725));
    equaln #(12) e2726(.a(buffered_input), .b(12'b101010100110), .eq(weq2726));
    equaln #(12) e2727(.a(buffered_input), .b(12'b101010100111), .eq(weq2727));
    equaln #(12) e2728(.a(buffered_input), .b(12'b101010101000), .eq(weq2728));
    equaln #(12) e2729(.a(buffered_input), .b(12'b101010101001), .eq(weq2729));
    equaln #(12) e2730(.a(buffered_input), .b(12'b101010101010), .eq(weq2730));
    equaln #(12) e2731(.a(buffered_input), .b(12'b101010101011), .eq(weq2731));
    equaln #(12) e2732(.a(buffered_input), .b(12'b101010101100), .eq(weq2732));
    equaln #(12) e2733(.a(buffered_input), .b(12'b101010101101), .eq(weq2733));
    equaln #(12) e2734(.a(buffered_input), .b(12'b101010101110), .eq(weq2734));
    equaln #(12) e2735(.a(buffered_input), .b(12'b101010101111), .eq(weq2735));
    equaln #(12) e2736(.a(buffered_input), .b(12'b101010110000), .eq(weq2736));
    equaln #(12) e2737(.a(buffered_input), .b(12'b101010110001), .eq(weq2737));
    equaln #(12) e2738(.a(buffered_input), .b(12'b101010110010), .eq(weq2738));
    equaln #(12) e2739(.a(buffered_input), .b(12'b101010110011), .eq(weq2739));
    equaln #(12) e2740(.a(buffered_input), .b(12'b101010110100), .eq(weq2740));
    equaln #(12) e2741(.a(buffered_input), .b(12'b101010110101), .eq(weq2741));
    equaln #(12) e2742(.a(buffered_input), .b(12'b101010110110), .eq(weq2742));
    equaln #(12) e2743(.a(buffered_input), .b(12'b101010110111), .eq(weq2743));
    equaln #(12) e2744(.a(buffered_input), .b(12'b101010111000), .eq(weq2744));
    equaln #(12) e2745(.a(buffered_input), .b(12'b101010111001), .eq(weq2745));
    equaln #(12) e2746(.a(buffered_input), .b(12'b101010111010), .eq(weq2746));
    equaln #(12) e2747(.a(buffered_input), .b(12'b101010111011), .eq(weq2747));
    equaln #(12) e2748(.a(buffered_input), .b(12'b101010111100), .eq(weq2748));
    equaln #(12) e2749(.a(buffered_input), .b(12'b101010111101), .eq(weq2749));
    equaln #(12) e2750(.a(buffered_input), .b(12'b101010111110), .eq(weq2750));
    equaln #(12) e2751(.a(buffered_input), .b(12'b101010111111), .eq(weq2751));
    equaln #(12) e2752(.a(buffered_input), .b(12'b101011000000), .eq(weq2752));
    equaln #(12) e2753(.a(buffered_input), .b(12'b101011000001), .eq(weq2753));
    equaln #(12) e2754(.a(buffered_input), .b(12'b101011000010), .eq(weq2754));
    equaln #(12) e2755(.a(buffered_input), .b(12'b101011000011), .eq(weq2755));
    equaln #(12) e2756(.a(buffered_input), .b(12'b101011000100), .eq(weq2756));
    equaln #(12) e2757(.a(buffered_input), .b(12'b101011000101), .eq(weq2757));
    equaln #(12) e2758(.a(buffered_input), .b(12'b101011000110), .eq(weq2758));
    equaln #(12) e2759(.a(buffered_input), .b(12'b101011000111), .eq(weq2759));
    equaln #(12) e2760(.a(buffered_input), .b(12'b101011001000), .eq(weq2760));
    equaln #(12) e2761(.a(buffered_input), .b(12'b101011001001), .eq(weq2761));
    equaln #(12) e2762(.a(buffered_input), .b(12'b101011001010), .eq(weq2762));
    equaln #(12) e2763(.a(buffered_input), .b(12'b101011001011), .eq(weq2763));
    equaln #(12) e2764(.a(buffered_input), .b(12'b101011001100), .eq(weq2764));
    equaln #(12) e2765(.a(buffered_input), .b(12'b101011001101), .eq(weq2765));
    equaln #(12) e2766(.a(buffered_input), .b(12'b101011001110), .eq(weq2766));
    equaln #(12) e2767(.a(buffered_input), .b(12'b101011001111), .eq(weq2767));
    equaln #(12) e2768(.a(buffered_input), .b(12'b101011010000), .eq(weq2768));
    equaln #(12) e2769(.a(buffered_input), .b(12'b101011010001), .eq(weq2769));
    equaln #(12) e2770(.a(buffered_input), .b(12'b101011010010), .eq(weq2770));
    equaln #(12) e2771(.a(buffered_input), .b(12'b101011010011), .eq(weq2771));
    equaln #(12) e2772(.a(buffered_input), .b(12'b101011010100), .eq(weq2772));
    equaln #(12) e2773(.a(buffered_input), .b(12'b101011010101), .eq(weq2773));
    equaln #(12) e2774(.a(buffered_input), .b(12'b101011010110), .eq(weq2774));
    equaln #(12) e2775(.a(buffered_input), .b(12'b101011010111), .eq(weq2775));
    equaln #(12) e2776(.a(buffered_input), .b(12'b101011011000), .eq(weq2776));
    equaln #(12) e2777(.a(buffered_input), .b(12'b101011011001), .eq(weq2777));
    equaln #(12) e2778(.a(buffered_input), .b(12'b101011011010), .eq(weq2778));
    equaln #(12) e2779(.a(buffered_input), .b(12'b101011011011), .eq(weq2779));
    equaln #(12) e2780(.a(buffered_input), .b(12'b101011011100), .eq(weq2780));
    equaln #(12) e2781(.a(buffered_input), .b(12'b101011011101), .eq(weq2781));
    equaln #(12) e2782(.a(buffered_input), .b(12'b101011011110), .eq(weq2782));
    equaln #(12) e2783(.a(buffered_input), .b(12'b101011011111), .eq(weq2783));
    equaln #(12) e2784(.a(buffered_input), .b(12'b101011100000), .eq(weq2784));
    equaln #(12) e2785(.a(buffered_input), .b(12'b101011100001), .eq(weq2785));
    equaln #(12) e2786(.a(buffered_input), .b(12'b101011100010), .eq(weq2786));
    equaln #(12) e2787(.a(buffered_input), .b(12'b101011100011), .eq(weq2787));
    equaln #(12) e2788(.a(buffered_input), .b(12'b101011100100), .eq(weq2788));
    equaln #(12) e2789(.a(buffered_input), .b(12'b101011100101), .eq(weq2789));
    equaln #(12) e2790(.a(buffered_input), .b(12'b101011100110), .eq(weq2790));
    equaln #(12) e2791(.a(buffered_input), .b(12'b101011100111), .eq(weq2791));
    equaln #(12) e2792(.a(buffered_input), .b(12'b101011101000), .eq(weq2792));
    equaln #(12) e2793(.a(buffered_input), .b(12'b101011101001), .eq(weq2793));
    equaln #(12) e2794(.a(buffered_input), .b(12'b101011101010), .eq(weq2794));
    equaln #(12) e2795(.a(buffered_input), .b(12'b101011101011), .eq(weq2795));
    equaln #(12) e2796(.a(buffered_input), .b(12'b101011101100), .eq(weq2796));
    equaln #(12) e2797(.a(buffered_input), .b(12'b101011101101), .eq(weq2797));
    equaln #(12) e2798(.a(buffered_input), .b(12'b101011101110), .eq(weq2798));
    equaln #(12) e2799(.a(buffered_input), .b(12'b101011101111), .eq(weq2799));
    equaln #(12) e2800(.a(buffered_input), .b(12'b101011110000), .eq(weq2800));
    equaln #(12) e2801(.a(buffered_input), .b(12'b101011110001), .eq(weq2801));
    equaln #(12) e2802(.a(buffered_input), .b(12'b101011110010), .eq(weq2802));
    equaln #(12) e2803(.a(buffered_input), .b(12'b101011110011), .eq(weq2803));
    equaln #(12) e2804(.a(buffered_input), .b(12'b101011110100), .eq(weq2804));
    equaln #(12) e2805(.a(buffered_input), .b(12'b101011110101), .eq(weq2805));
    equaln #(12) e2806(.a(buffered_input), .b(12'b101011110110), .eq(weq2806));
    equaln #(12) e2807(.a(buffered_input), .b(12'b101011110111), .eq(weq2807));
    equaln #(12) e2808(.a(buffered_input), .b(12'b101011111000), .eq(weq2808));
    equaln #(12) e2809(.a(buffered_input), .b(12'b101011111001), .eq(weq2809));
    equaln #(12) e2810(.a(buffered_input), .b(12'b101011111010), .eq(weq2810));
    equaln #(12) e2811(.a(buffered_input), .b(12'b101011111011), .eq(weq2811));
    equaln #(12) e2812(.a(buffered_input), .b(12'b101011111100), .eq(weq2812));
    equaln #(12) e2813(.a(buffered_input), .b(12'b101011111101), .eq(weq2813));
    equaln #(12) e2814(.a(buffered_input), .b(12'b101011111110), .eq(weq2814));
    equaln #(12) e2815(.a(buffered_input), .b(12'b101011111111), .eq(weq2815));
    equaln #(12) e2816(.a(buffered_input), .b(12'b101100000000), .eq(weq2816));
    equaln #(12) e2817(.a(buffered_input), .b(12'b101100000001), .eq(weq2817));
    equaln #(12) e2818(.a(buffered_input), .b(12'b101100000010), .eq(weq2818));
    equaln #(12) e2819(.a(buffered_input), .b(12'b101100000011), .eq(weq2819));
    equaln #(12) e2820(.a(buffered_input), .b(12'b101100000100), .eq(weq2820));
    equaln #(12) e2821(.a(buffered_input), .b(12'b101100000101), .eq(weq2821));
    equaln #(12) e2822(.a(buffered_input), .b(12'b101100000110), .eq(weq2822));
    equaln #(12) e2823(.a(buffered_input), .b(12'b101100000111), .eq(weq2823));
    equaln #(12) e2824(.a(buffered_input), .b(12'b101100001000), .eq(weq2824));
    equaln #(12) e2825(.a(buffered_input), .b(12'b101100001001), .eq(weq2825));
    equaln #(12) e2826(.a(buffered_input), .b(12'b101100001010), .eq(weq2826));
    equaln #(12) e2827(.a(buffered_input), .b(12'b101100001011), .eq(weq2827));
    equaln #(12) e2828(.a(buffered_input), .b(12'b101100001100), .eq(weq2828));
    equaln #(12) e2829(.a(buffered_input), .b(12'b101100001101), .eq(weq2829));
    equaln #(12) e2830(.a(buffered_input), .b(12'b101100001110), .eq(weq2830));
    equaln #(12) e2831(.a(buffered_input), .b(12'b101100001111), .eq(weq2831));
    equaln #(12) e2832(.a(buffered_input), .b(12'b101100010000), .eq(weq2832));
    equaln #(12) e2833(.a(buffered_input), .b(12'b101100010001), .eq(weq2833));
    equaln #(12) e2834(.a(buffered_input), .b(12'b101100010010), .eq(weq2834));
    equaln #(12) e2835(.a(buffered_input), .b(12'b101100010011), .eq(weq2835));
    equaln #(12) e2836(.a(buffered_input), .b(12'b101100010100), .eq(weq2836));
    equaln #(12) e2837(.a(buffered_input), .b(12'b101100010101), .eq(weq2837));
    equaln #(12) e2838(.a(buffered_input), .b(12'b101100010110), .eq(weq2838));
    equaln #(12) e2839(.a(buffered_input), .b(12'b101100010111), .eq(weq2839));
    equaln #(12) e2840(.a(buffered_input), .b(12'b101100011000), .eq(weq2840));
    equaln #(12) e2841(.a(buffered_input), .b(12'b101100011001), .eq(weq2841));
    equaln #(12) e2842(.a(buffered_input), .b(12'b101100011010), .eq(weq2842));
    equaln #(12) e2843(.a(buffered_input), .b(12'b101100011011), .eq(weq2843));
    equaln #(12) e2844(.a(buffered_input), .b(12'b101100011100), .eq(weq2844));
    equaln #(12) e2845(.a(buffered_input), .b(12'b101100011101), .eq(weq2845));
    equaln #(12) e2846(.a(buffered_input), .b(12'b101100011110), .eq(weq2846));
    equaln #(12) e2847(.a(buffered_input), .b(12'b101100011111), .eq(weq2847));
    equaln #(12) e2848(.a(buffered_input), .b(12'b101100100000), .eq(weq2848));
    equaln #(12) e2849(.a(buffered_input), .b(12'b101100100001), .eq(weq2849));
    equaln #(12) e2850(.a(buffered_input), .b(12'b101100100010), .eq(weq2850));
    equaln #(12) e2851(.a(buffered_input), .b(12'b101100100011), .eq(weq2851));
    equaln #(12) e2852(.a(buffered_input), .b(12'b101100100100), .eq(weq2852));
    equaln #(12) e2853(.a(buffered_input), .b(12'b101100100101), .eq(weq2853));
    equaln #(12) e2854(.a(buffered_input), .b(12'b101100100110), .eq(weq2854));
    equaln #(12) e2855(.a(buffered_input), .b(12'b101100100111), .eq(weq2855));
    equaln #(12) e2856(.a(buffered_input), .b(12'b101100101000), .eq(weq2856));
    equaln #(12) e2857(.a(buffered_input), .b(12'b101100101001), .eq(weq2857));
    equaln #(12) e2858(.a(buffered_input), .b(12'b101100101010), .eq(weq2858));
    equaln #(12) e2859(.a(buffered_input), .b(12'b101100101011), .eq(weq2859));
    equaln #(12) e2860(.a(buffered_input), .b(12'b101100101100), .eq(weq2860));
    equaln #(12) e2861(.a(buffered_input), .b(12'b101100101101), .eq(weq2861));
    equaln #(12) e2862(.a(buffered_input), .b(12'b101100101110), .eq(weq2862));
    equaln #(12) e2863(.a(buffered_input), .b(12'b101100101111), .eq(weq2863));
    equaln #(12) e2864(.a(buffered_input), .b(12'b101100110000), .eq(weq2864));
    equaln #(12) e2865(.a(buffered_input), .b(12'b101100110001), .eq(weq2865));
    equaln #(12) e2866(.a(buffered_input), .b(12'b101100110010), .eq(weq2866));
    equaln #(12) e2867(.a(buffered_input), .b(12'b101100110011), .eq(weq2867));
    equaln #(12) e2868(.a(buffered_input), .b(12'b101100110100), .eq(weq2868));
    equaln #(12) e2869(.a(buffered_input), .b(12'b101100110101), .eq(weq2869));
    equaln #(12) e2870(.a(buffered_input), .b(12'b101100110110), .eq(weq2870));
    equaln #(12) e2871(.a(buffered_input), .b(12'b101100110111), .eq(weq2871));
    equaln #(12) e2872(.a(buffered_input), .b(12'b101100111000), .eq(weq2872));
    equaln #(12) e2873(.a(buffered_input), .b(12'b101100111001), .eq(weq2873));
    equaln #(12) e2874(.a(buffered_input), .b(12'b101100111010), .eq(weq2874));
    equaln #(12) e2875(.a(buffered_input), .b(12'b101100111011), .eq(weq2875));
    equaln #(12) e2876(.a(buffered_input), .b(12'b101100111100), .eq(weq2876));
    equaln #(12) e2877(.a(buffered_input), .b(12'b101100111101), .eq(weq2877));
    equaln #(12) e2878(.a(buffered_input), .b(12'b101100111110), .eq(weq2878));
    equaln #(12) e2879(.a(buffered_input), .b(12'b101100111111), .eq(weq2879));
    equaln #(12) e2880(.a(buffered_input), .b(12'b101101000000), .eq(weq2880));
    equaln #(12) e2881(.a(buffered_input), .b(12'b101101000001), .eq(weq2881));
    equaln #(12) e2882(.a(buffered_input), .b(12'b101101000010), .eq(weq2882));
    equaln #(12) e2883(.a(buffered_input), .b(12'b101101000011), .eq(weq2883));
    equaln #(12) e2884(.a(buffered_input), .b(12'b101101000100), .eq(weq2884));
    equaln #(12) e2885(.a(buffered_input), .b(12'b101101000101), .eq(weq2885));
    equaln #(12) e2886(.a(buffered_input), .b(12'b101101000110), .eq(weq2886));
    equaln #(12) e2887(.a(buffered_input), .b(12'b101101000111), .eq(weq2887));
    equaln #(12) e2888(.a(buffered_input), .b(12'b101101001000), .eq(weq2888));
    equaln #(12) e2889(.a(buffered_input), .b(12'b101101001001), .eq(weq2889));
    equaln #(12) e2890(.a(buffered_input), .b(12'b101101001010), .eq(weq2890));
    equaln #(12) e2891(.a(buffered_input), .b(12'b101101001011), .eq(weq2891));
    equaln #(12) e2892(.a(buffered_input), .b(12'b101101001100), .eq(weq2892));
    equaln #(12) e2893(.a(buffered_input), .b(12'b101101001101), .eq(weq2893));
    equaln #(12) e2894(.a(buffered_input), .b(12'b101101001110), .eq(weq2894));
    equaln #(12) e2895(.a(buffered_input), .b(12'b101101001111), .eq(weq2895));
    equaln #(12) e2896(.a(buffered_input), .b(12'b101101010000), .eq(weq2896));
    equaln #(12) e2897(.a(buffered_input), .b(12'b101101010001), .eq(weq2897));
    equaln #(12) e2898(.a(buffered_input), .b(12'b101101010010), .eq(weq2898));
    equaln #(12) e2899(.a(buffered_input), .b(12'b101101010011), .eq(weq2899));
    equaln #(12) e2900(.a(buffered_input), .b(12'b101101010100), .eq(weq2900));
    equaln #(12) e2901(.a(buffered_input), .b(12'b101101010101), .eq(weq2901));
    equaln #(12) e2902(.a(buffered_input), .b(12'b101101010110), .eq(weq2902));
    equaln #(12) e2903(.a(buffered_input), .b(12'b101101010111), .eq(weq2903));
    equaln #(12) e2904(.a(buffered_input), .b(12'b101101011000), .eq(weq2904));
    equaln #(12) e2905(.a(buffered_input), .b(12'b101101011001), .eq(weq2905));
    equaln #(12) e2906(.a(buffered_input), .b(12'b101101011010), .eq(weq2906));
    equaln #(12) e2907(.a(buffered_input), .b(12'b101101011011), .eq(weq2907));
    equaln #(12) e2908(.a(buffered_input), .b(12'b101101011100), .eq(weq2908));
    equaln #(12) e2909(.a(buffered_input), .b(12'b101101011101), .eq(weq2909));
    equaln #(12) e2910(.a(buffered_input), .b(12'b101101011110), .eq(weq2910));
    equaln #(12) e2911(.a(buffered_input), .b(12'b101101011111), .eq(weq2911));
    equaln #(12) e2912(.a(buffered_input), .b(12'b101101100000), .eq(weq2912));
    equaln #(12) e2913(.a(buffered_input), .b(12'b101101100001), .eq(weq2913));
    equaln #(12) e2914(.a(buffered_input), .b(12'b101101100010), .eq(weq2914));
    equaln #(12) e2915(.a(buffered_input), .b(12'b101101100011), .eq(weq2915));
    equaln #(12) e2916(.a(buffered_input), .b(12'b101101100100), .eq(weq2916));
    equaln #(12) e2917(.a(buffered_input), .b(12'b101101100101), .eq(weq2917));
    equaln #(12) e2918(.a(buffered_input), .b(12'b101101100110), .eq(weq2918));
    equaln #(12) e2919(.a(buffered_input), .b(12'b101101100111), .eq(weq2919));
    equaln #(12) e2920(.a(buffered_input), .b(12'b101101101000), .eq(weq2920));
    equaln #(12) e2921(.a(buffered_input), .b(12'b101101101001), .eq(weq2921));
    equaln #(12) e2922(.a(buffered_input), .b(12'b101101101010), .eq(weq2922));
    equaln #(12) e2923(.a(buffered_input), .b(12'b101101101011), .eq(weq2923));
    equaln #(12) e2924(.a(buffered_input), .b(12'b101101101100), .eq(weq2924));
    equaln #(12) e2925(.a(buffered_input), .b(12'b101101101101), .eq(weq2925));
    equaln #(12) e2926(.a(buffered_input), .b(12'b101101101110), .eq(weq2926));
    equaln #(12) e2927(.a(buffered_input), .b(12'b101101101111), .eq(weq2927));
    equaln #(12) e2928(.a(buffered_input), .b(12'b101101110000), .eq(weq2928));
    equaln #(12) e2929(.a(buffered_input), .b(12'b101101110001), .eq(weq2929));
    equaln #(12) e2930(.a(buffered_input), .b(12'b101101110010), .eq(weq2930));
    equaln #(12) e2931(.a(buffered_input), .b(12'b101101110011), .eq(weq2931));
    equaln #(12) e2932(.a(buffered_input), .b(12'b101101110100), .eq(weq2932));
    equaln #(12) e2933(.a(buffered_input), .b(12'b101101110101), .eq(weq2933));
    equaln #(12) e2934(.a(buffered_input), .b(12'b101101110110), .eq(weq2934));
    equaln #(12) e2935(.a(buffered_input), .b(12'b101101110111), .eq(weq2935));
    equaln #(12) e2936(.a(buffered_input), .b(12'b101101111000), .eq(weq2936));
    equaln #(12) e2937(.a(buffered_input), .b(12'b101101111001), .eq(weq2937));
    equaln #(12) e2938(.a(buffered_input), .b(12'b101101111010), .eq(weq2938));
    equaln #(12) e2939(.a(buffered_input), .b(12'b101101111011), .eq(weq2939));
    equaln #(12) e2940(.a(buffered_input), .b(12'b101101111100), .eq(weq2940));
    equaln #(12) e2941(.a(buffered_input), .b(12'b101101111101), .eq(weq2941));
    equaln #(12) e2942(.a(buffered_input), .b(12'b101101111110), .eq(weq2942));
    equaln #(12) e2943(.a(buffered_input), .b(12'b101101111111), .eq(weq2943));
    equaln #(12) e2944(.a(buffered_input), .b(12'b101110000000), .eq(weq2944));
    equaln #(12) e2945(.a(buffered_input), .b(12'b101110000001), .eq(weq2945));
    equaln #(12) e2946(.a(buffered_input), .b(12'b101110000010), .eq(weq2946));
    equaln #(12) e2947(.a(buffered_input), .b(12'b101110000011), .eq(weq2947));
    equaln #(12) e2948(.a(buffered_input), .b(12'b101110000100), .eq(weq2948));
    equaln #(12) e2949(.a(buffered_input), .b(12'b101110000101), .eq(weq2949));
    equaln #(12) e2950(.a(buffered_input), .b(12'b101110000110), .eq(weq2950));
    equaln #(12) e2951(.a(buffered_input), .b(12'b101110000111), .eq(weq2951));
    equaln #(12) e2952(.a(buffered_input), .b(12'b101110001000), .eq(weq2952));
    equaln #(12) e2953(.a(buffered_input), .b(12'b101110001001), .eq(weq2953));
    equaln #(12) e2954(.a(buffered_input), .b(12'b101110001010), .eq(weq2954));
    equaln #(12) e2955(.a(buffered_input), .b(12'b101110001011), .eq(weq2955));
    equaln #(12) e2956(.a(buffered_input), .b(12'b101110001100), .eq(weq2956));
    equaln #(12) e2957(.a(buffered_input), .b(12'b101110001101), .eq(weq2957));
    equaln #(12) e2958(.a(buffered_input), .b(12'b101110001110), .eq(weq2958));
    equaln #(12) e2959(.a(buffered_input), .b(12'b101110001111), .eq(weq2959));
    equaln #(12) e2960(.a(buffered_input), .b(12'b101110010000), .eq(weq2960));
    equaln #(12) e2961(.a(buffered_input), .b(12'b101110010001), .eq(weq2961));
    equaln #(12) e2962(.a(buffered_input), .b(12'b101110010010), .eq(weq2962));
    equaln #(12) e2963(.a(buffered_input), .b(12'b101110010011), .eq(weq2963));
    equaln #(12) e2964(.a(buffered_input), .b(12'b101110010100), .eq(weq2964));
    equaln #(12) e2965(.a(buffered_input), .b(12'b101110010101), .eq(weq2965));
    equaln #(12) e2966(.a(buffered_input), .b(12'b101110010110), .eq(weq2966));
    equaln #(12) e2967(.a(buffered_input), .b(12'b101110010111), .eq(weq2967));
    equaln #(12) e2968(.a(buffered_input), .b(12'b101110011000), .eq(weq2968));
    equaln #(12) e2969(.a(buffered_input), .b(12'b101110011001), .eq(weq2969));
    equaln #(12) e2970(.a(buffered_input), .b(12'b101110011010), .eq(weq2970));
    equaln #(12) e2971(.a(buffered_input), .b(12'b101110011011), .eq(weq2971));
    equaln #(12) e2972(.a(buffered_input), .b(12'b101110011100), .eq(weq2972));
    equaln #(12) e2973(.a(buffered_input), .b(12'b101110011101), .eq(weq2973));
    equaln #(12) e2974(.a(buffered_input), .b(12'b101110011110), .eq(weq2974));
    equaln #(12) e2975(.a(buffered_input), .b(12'b101110011111), .eq(weq2975));
    equaln #(12) e2976(.a(buffered_input), .b(12'b101110100000), .eq(weq2976));
    equaln #(12) e2977(.a(buffered_input), .b(12'b101110100001), .eq(weq2977));
    equaln #(12) e2978(.a(buffered_input), .b(12'b101110100010), .eq(weq2978));
    equaln #(12) e2979(.a(buffered_input), .b(12'b101110100011), .eq(weq2979));
    equaln #(12) e2980(.a(buffered_input), .b(12'b101110100100), .eq(weq2980));
    equaln #(12) e2981(.a(buffered_input), .b(12'b101110100101), .eq(weq2981));
    equaln #(12) e2982(.a(buffered_input), .b(12'b101110100110), .eq(weq2982));
    equaln #(12) e2983(.a(buffered_input), .b(12'b101110100111), .eq(weq2983));
    equaln #(12) e2984(.a(buffered_input), .b(12'b101110101000), .eq(weq2984));
    equaln #(12) e2985(.a(buffered_input), .b(12'b101110101001), .eq(weq2985));
    equaln #(12) e2986(.a(buffered_input), .b(12'b101110101010), .eq(weq2986));
    equaln #(12) e2987(.a(buffered_input), .b(12'b101110101011), .eq(weq2987));
    equaln #(12) e2988(.a(buffered_input), .b(12'b101110101100), .eq(weq2988));
    equaln #(12) e2989(.a(buffered_input), .b(12'b101110101101), .eq(weq2989));
    equaln #(12) e2990(.a(buffered_input), .b(12'b101110101110), .eq(weq2990));
    equaln #(12) e2991(.a(buffered_input), .b(12'b101110101111), .eq(weq2991));
    equaln #(12) e2992(.a(buffered_input), .b(12'b101110110000), .eq(weq2992));
    equaln #(12) e2993(.a(buffered_input), .b(12'b101110110001), .eq(weq2993));
    equaln #(12) e2994(.a(buffered_input), .b(12'b101110110010), .eq(weq2994));
    equaln #(12) e2995(.a(buffered_input), .b(12'b101110110011), .eq(weq2995));
    equaln #(12) e2996(.a(buffered_input), .b(12'b101110110100), .eq(weq2996));
    equaln #(12) e2997(.a(buffered_input), .b(12'b101110110101), .eq(weq2997));
    equaln #(12) e2998(.a(buffered_input), .b(12'b101110110110), .eq(weq2998));
    equaln #(12) e2999(.a(buffered_input), .b(12'b101110110111), .eq(weq2999));
    equaln #(12) e3000(.a(buffered_input), .b(12'b101110111000), .eq(weq3000));
    equaln #(12) e3001(.a(buffered_input), .b(12'b101110111001), .eq(weq3001));
    equaln #(12) e3002(.a(buffered_input), .b(12'b101110111010), .eq(weq3002));
    equaln #(12) e3003(.a(buffered_input), .b(12'b101110111011), .eq(weq3003));
    equaln #(12) e3004(.a(buffered_input), .b(12'b101110111100), .eq(weq3004));
    equaln #(12) e3005(.a(buffered_input), .b(12'b101110111101), .eq(weq3005));
    equaln #(12) e3006(.a(buffered_input), .b(12'b101110111110), .eq(weq3006));
    equaln #(12) e3007(.a(buffered_input), .b(12'b101110111111), .eq(weq3007));
    equaln #(12) e3008(.a(buffered_input), .b(12'b101111000000), .eq(weq3008));
    equaln #(12) e3009(.a(buffered_input), .b(12'b101111000001), .eq(weq3009));
    equaln #(12) e3010(.a(buffered_input), .b(12'b101111000010), .eq(weq3010));
    equaln #(12) e3011(.a(buffered_input), .b(12'b101111000011), .eq(weq3011));
    equaln #(12) e3012(.a(buffered_input), .b(12'b101111000100), .eq(weq3012));
    equaln #(12) e3013(.a(buffered_input), .b(12'b101111000101), .eq(weq3013));
    equaln #(12) e3014(.a(buffered_input), .b(12'b101111000110), .eq(weq3014));
    equaln #(12) e3015(.a(buffered_input), .b(12'b101111000111), .eq(weq3015));
    equaln #(12) e3016(.a(buffered_input), .b(12'b101111001000), .eq(weq3016));
    equaln #(12) e3017(.a(buffered_input), .b(12'b101111001001), .eq(weq3017));
    equaln #(12) e3018(.a(buffered_input), .b(12'b101111001010), .eq(weq3018));
    equaln #(12) e3019(.a(buffered_input), .b(12'b101111001011), .eq(weq3019));
    equaln #(12) e3020(.a(buffered_input), .b(12'b101111001100), .eq(weq3020));
    equaln #(12) e3021(.a(buffered_input), .b(12'b101111001101), .eq(weq3021));
    equaln #(12) e3022(.a(buffered_input), .b(12'b101111001110), .eq(weq3022));
    equaln #(12) e3023(.a(buffered_input), .b(12'b101111001111), .eq(weq3023));
    equaln #(12) e3024(.a(buffered_input), .b(12'b101111010000), .eq(weq3024));
    equaln #(12) e3025(.a(buffered_input), .b(12'b101111010001), .eq(weq3025));
    equaln #(12) e3026(.a(buffered_input), .b(12'b101111010010), .eq(weq3026));
    equaln #(12) e3027(.a(buffered_input), .b(12'b101111010011), .eq(weq3027));
    equaln #(12) e3028(.a(buffered_input), .b(12'b101111010100), .eq(weq3028));
    equaln #(12) e3029(.a(buffered_input), .b(12'b101111010101), .eq(weq3029));
    equaln #(12) e3030(.a(buffered_input), .b(12'b101111010110), .eq(weq3030));
    equaln #(12) e3031(.a(buffered_input), .b(12'b101111010111), .eq(weq3031));
    equaln #(12) e3032(.a(buffered_input), .b(12'b101111011000), .eq(weq3032));
    equaln #(12) e3033(.a(buffered_input), .b(12'b101111011001), .eq(weq3033));
    equaln #(12) e3034(.a(buffered_input), .b(12'b101111011010), .eq(weq3034));
    equaln #(12) e3035(.a(buffered_input), .b(12'b101111011011), .eq(weq3035));
    equaln #(12) e3036(.a(buffered_input), .b(12'b101111011100), .eq(weq3036));
    equaln #(12) e3037(.a(buffered_input), .b(12'b101111011101), .eq(weq3037));
    equaln #(12) e3038(.a(buffered_input), .b(12'b101111011110), .eq(weq3038));
    equaln #(12) e3039(.a(buffered_input), .b(12'b101111011111), .eq(weq3039));
    equaln #(12) e3040(.a(buffered_input), .b(12'b101111100000), .eq(weq3040));
    equaln #(12) e3041(.a(buffered_input), .b(12'b101111100001), .eq(weq3041));
    equaln #(12) e3042(.a(buffered_input), .b(12'b101111100010), .eq(weq3042));
    equaln #(12) e3043(.a(buffered_input), .b(12'b101111100011), .eq(weq3043));
    equaln #(12) e3044(.a(buffered_input), .b(12'b101111100100), .eq(weq3044));
    equaln #(12) e3045(.a(buffered_input), .b(12'b101111100101), .eq(weq3045));
    equaln #(12) e3046(.a(buffered_input), .b(12'b101111100110), .eq(weq3046));
    equaln #(12) e3047(.a(buffered_input), .b(12'b101111100111), .eq(weq3047));
    equaln #(12) e3048(.a(buffered_input), .b(12'b101111101000), .eq(weq3048));
    equaln #(12) e3049(.a(buffered_input), .b(12'b101111101001), .eq(weq3049));
    equaln #(12) e3050(.a(buffered_input), .b(12'b101111101010), .eq(weq3050));
    equaln #(12) e3051(.a(buffered_input), .b(12'b101111101011), .eq(weq3051));
    equaln #(12) e3052(.a(buffered_input), .b(12'b101111101100), .eq(weq3052));
    equaln #(12) e3053(.a(buffered_input), .b(12'b101111101101), .eq(weq3053));
    equaln #(12) e3054(.a(buffered_input), .b(12'b101111101110), .eq(weq3054));
    equaln #(12) e3055(.a(buffered_input), .b(12'b101111101111), .eq(weq3055));
    equaln #(12) e3056(.a(buffered_input), .b(12'b101111110000), .eq(weq3056));
    equaln #(12) e3057(.a(buffered_input), .b(12'b101111110001), .eq(weq3057));
    equaln #(12) e3058(.a(buffered_input), .b(12'b101111110010), .eq(weq3058));
    equaln #(12) e3059(.a(buffered_input), .b(12'b101111110011), .eq(weq3059));
    equaln #(12) e3060(.a(buffered_input), .b(12'b101111110100), .eq(weq3060));
    equaln #(12) e3061(.a(buffered_input), .b(12'b101111110101), .eq(weq3061));
    equaln #(12) e3062(.a(buffered_input), .b(12'b101111110110), .eq(weq3062));
    equaln #(12) e3063(.a(buffered_input), .b(12'b101111110111), .eq(weq3063));
    equaln #(12) e3064(.a(buffered_input), .b(12'b101111111000), .eq(weq3064));
    equaln #(12) e3065(.a(buffered_input), .b(12'b101111111001), .eq(weq3065));
    equaln #(12) e3066(.a(buffered_input), .b(12'b101111111010), .eq(weq3066));
    equaln #(12) e3067(.a(buffered_input), .b(12'b101111111011), .eq(weq3067));
    equaln #(12) e3068(.a(buffered_input), .b(12'b101111111100), .eq(weq3068));
    equaln #(12) e3069(.a(buffered_input), .b(12'b101111111101), .eq(weq3069));
    equaln #(12) e3070(.a(buffered_input), .b(12'b101111111110), .eq(weq3070));
    equaln #(12) e3071(.a(buffered_input), .b(12'b101111111111), .eq(weq3071));
    equaln #(12) e3072(.a(buffered_input), .b(12'b110000000000), .eq(weq3072));
    equaln #(12) e3073(.a(buffered_input), .b(12'b110000000001), .eq(weq3073));
    equaln #(12) e3074(.a(buffered_input), .b(12'b110000000010), .eq(weq3074));
    equaln #(12) e3075(.a(buffered_input), .b(12'b110000000011), .eq(weq3075));
    equaln #(12) e3076(.a(buffered_input), .b(12'b110000000100), .eq(weq3076));
    equaln #(12) e3077(.a(buffered_input), .b(12'b110000000101), .eq(weq3077));
    equaln #(12) e3078(.a(buffered_input), .b(12'b110000000110), .eq(weq3078));
    equaln #(12) e3079(.a(buffered_input), .b(12'b110000000111), .eq(weq3079));
    equaln #(12) e3080(.a(buffered_input), .b(12'b110000001000), .eq(weq3080));
    equaln #(12) e3081(.a(buffered_input), .b(12'b110000001001), .eq(weq3081));
    equaln #(12) e3082(.a(buffered_input), .b(12'b110000001010), .eq(weq3082));
    equaln #(12) e3083(.a(buffered_input), .b(12'b110000001011), .eq(weq3083));
    equaln #(12) e3084(.a(buffered_input), .b(12'b110000001100), .eq(weq3084));
    equaln #(12) e3085(.a(buffered_input), .b(12'b110000001101), .eq(weq3085));
    equaln #(12) e3086(.a(buffered_input), .b(12'b110000001110), .eq(weq3086));
    equaln #(12) e3087(.a(buffered_input), .b(12'b110000001111), .eq(weq3087));
    equaln #(12) e3088(.a(buffered_input), .b(12'b110000010000), .eq(weq3088));
    equaln #(12) e3089(.a(buffered_input), .b(12'b110000010001), .eq(weq3089));
    equaln #(12) e3090(.a(buffered_input), .b(12'b110000010010), .eq(weq3090));
    equaln #(12) e3091(.a(buffered_input), .b(12'b110000010011), .eq(weq3091));
    equaln #(12) e3092(.a(buffered_input), .b(12'b110000010100), .eq(weq3092));
    equaln #(12) e3093(.a(buffered_input), .b(12'b110000010101), .eq(weq3093));
    equaln #(12) e3094(.a(buffered_input), .b(12'b110000010110), .eq(weq3094));
    equaln #(12) e3095(.a(buffered_input), .b(12'b110000010111), .eq(weq3095));
    equaln #(12) e3096(.a(buffered_input), .b(12'b110000011000), .eq(weq3096));
    equaln #(12) e3097(.a(buffered_input), .b(12'b110000011001), .eq(weq3097));
    equaln #(12) e3098(.a(buffered_input), .b(12'b110000011010), .eq(weq3098));
    equaln #(12) e3099(.a(buffered_input), .b(12'b110000011011), .eq(weq3099));
    equaln #(12) e3100(.a(buffered_input), .b(12'b110000011100), .eq(weq3100));
    equaln #(12) e3101(.a(buffered_input), .b(12'b110000011101), .eq(weq3101));
    equaln #(12) e3102(.a(buffered_input), .b(12'b110000011110), .eq(weq3102));
    equaln #(12) e3103(.a(buffered_input), .b(12'b110000011111), .eq(weq3103));
    equaln #(12) e3104(.a(buffered_input), .b(12'b110000100000), .eq(weq3104));
    equaln #(12) e3105(.a(buffered_input), .b(12'b110000100001), .eq(weq3105));
    equaln #(12) e3106(.a(buffered_input), .b(12'b110000100010), .eq(weq3106));
    equaln #(12) e3107(.a(buffered_input), .b(12'b110000100011), .eq(weq3107));
    equaln #(12) e3108(.a(buffered_input), .b(12'b110000100100), .eq(weq3108));
    equaln #(12) e3109(.a(buffered_input), .b(12'b110000100101), .eq(weq3109));
    equaln #(12) e3110(.a(buffered_input), .b(12'b110000100110), .eq(weq3110));
    equaln #(12) e3111(.a(buffered_input), .b(12'b110000100111), .eq(weq3111));
    equaln #(12) e3112(.a(buffered_input), .b(12'b110000101000), .eq(weq3112));
    equaln #(12) e3113(.a(buffered_input), .b(12'b110000101001), .eq(weq3113));
    equaln #(12) e3114(.a(buffered_input), .b(12'b110000101010), .eq(weq3114));
    equaln #(12) e3115(.a(buffered_input), .b(12'b110000101011), .eq(weq3115));
    equaln #(12) e3116(.a(buffered_input), .b(12'b110000101100), .eq(weq3116));
    equaln #(12) e3117(.a(buffered_input), .b(12'b110000101101), .eq(weq3117));
    equaln #(12) e3118(.a(buffered_input), .b(12'b110000101110), .eq(weq3118));
    equaln #(12) e3119(.a(buffered_input), .b(12'b110000101111), .eq(weq3119));
    equaln #(12) e3120(.a(buffered_input), .b(12'b110000110000), .eq(weq3120));
    equaln #(12) e3121(.a(buffered_input), .b(12'b110000110001), .eq(weq3121));
    equaln #(12) e3122(.a(buffered_input), .b(12'b110000110010), .eq(weq3122));
    equaln #(12) e3123(.a(buffered_input), .b(12'b110000110011), .eq(weq3123));
    equaln #(12) e3124(.a(buffered_input), .b(12'b110000110100), .eq(weq3124));
    equaln #(12) e3125(.a(buffered_input), .b(12'b110000110101), .eq(weq3125));
    equaln #(12) e3126(.a(buffered_input), .b(12'b110000110110), .eq(weq3126));
    equaln #(12) e3127(.a(buffered_input), .b(12'b110000110111), .eq(weq3127));
    equaln #(12) e3128(.a(buffered_input), .b(12'b110000111000), .eq(weq3128));
    equaln #(12) e3129(.a(buffered_input), .b(12'b110000111001), .eq(weq3129));
    equaln #(12) e3130(.a(buffered_input), .b(12'b110000111010), .eq(weq3130));
    equaln #(12) e3131(.a(buffered_input), .b(12'b110000111011), .eq(weq3131));
    equaln #(12) e3132(.a(buffered_input), .b(12'b110000111100), .eq(weq3132));
    equaln #(12) e3133(.a(buffered_input), .b(12'b110000111101), .eq(weq3133));
    equaln #(12) e3134(.a(buffered_input), .b(12'b110000111110), .eq(weq3134));
    equaln #(12) e3135(.a(buffered_input), .b(12'b110000111111), .eq(weq3135));
    equaln #(12) e3136(.a(buffered_input), .b(12'b110001000000), .eq(weq3136));
    equaln #(12) e3137(.a(buffered_input), .b(12'b110001000001), .eq(weq3137));
    equaln #(12) e3138(.a(buffered_input), .b(12'b110001000010), .eq(weq3138));
    equaln #(12) e3139(.a(buffered_input), .b(12'b110001000011), .eq(weq3139));
    equaln #(12) e3140(.a(buffered_input), .b(12'b110001000100), .eq(weq3140));
    equaln #(12) e3141(.a(buffered_input), .b(12'b110001000101), .eq(weq3141));
    equaln #(12) e3142(.a(buffered_input), .b(12'b110001000110), .eq(weq3142));
    equaln #(12) e3143(.a(buffered_input), .b(12'b110001000111), .eq(weq3143));
    equaln #(12) e3144(.a(buffered_input), .b(12'b110001001000), .eq(weq3144));
    equaln #(12) e3145(.a(buffered_input), .b(12'b110001001001), .eq(weq3145));
    equaln #(12) e3146(.a(buffered_input), .b(12'b110001001010), .eq(weq3146));
    equaln #(12) e3147(.a(buffered_input), .b(12'b110001001011), .eq(weq3147));
    equaln #(12) e3148(.a(buffered_input), .b(12'b110001001100), .eq(weq3148));
    equaln #(12) e3149(.a(buffered_input), .b(12'b110001001101), .eq(weq3149));
    equaln #(12) e3150(.a(buffered_input), .b(12'b110001001110), .eq(weq3150));
    equaln #(12) e3151(.a(buffered_input), .b(12'b110001001111), .eq(weq3151));
    equaln #(12) e3152(.a(buffered_input), .b(12'b110001010000), .eq(weq3152));
    equaln #(12) e3153(.a(buffered_input), .b(12'b110001010001), .eq(weq3153));
    equaln #(12) e3154(.a(buffered_input), .b(12'b110001010010), .eq(weq3154));
    equaln #(12) e3155(.a(buffered_input), .b(12'b110001010011), .eq(weq3155));
    equaln #(12) e3156(.a(buffered_input), .b(12'b110001010100), .eq(weq3156));
    equaln #(12) e3157(.a(buffered_input), .b(12'b110001010101), .eq(weq3157));
    equaln #(12) e3158(.a(buffered_input), .b(12'b110001010110), .eq(weq3158));
    equaln #(12) e3159(.a(buffered_input), .b(12'b110001010111), .eq(weq3159));
    equaln #(12) e3160(.a(buffered_input), .b(12'b110001011000), .eq(weq3160));
    equaln #(12) e3161(.a(buffered_input), .b(12'b110001011001), .eq(weq3161));
    equaln #(12) e3162(.a(buffered_input), .b(12'b110001011010), .eq(weq3162));
    equaln #(12) e3163(.a(buffered_input), .b(12'b110001011011), .eq(weq3163));
    equaln #(12) e3164(.a(buffered_input), .b(12'b110001011100), .eq(weq3164));
    equaln #(12) e3165(.a(buffered_input), .b(12'b110001011101), .eq(weq3165));
    equaln #(12) e3166(.a(buffered_input), .b(12'b110001011110), .eq(weq3166));
    equaln #(12) e3167(.a(buffered_input), .b(12'b110001011111), .eq(weq3167));
    equaln #(12) e3168(.a(buffered_input), .b(12'b110001100000), .eq(weq3168));
    equaln #(12) e3169(.a(buffered_input), .b(12'b110001100001), .eq(weq3169));
    equaln #(12) e3170(.a(buffered_input), .b(12'b110001100010), .eq(weq3170));
    equaln #(12) e3171(.a(buffered_input), .b(12'b110001100011), .eq(weq3171));
    equaln #(12) e3172(.a(buffered_input), .b(12'b110001100100), .eq(weq3172));
    equaln #(12) e3173(.a(buffered_input), .b(12'b110001100101), .eq(weq3173));
    equaln #(12) e3174(.a(buffered_input), .b(12'b110001100110), .eq(weq3174));
    equaln #(12) e3175(.a(buffered_input), .b(12'b110001100111), .eq(weq3175));
    equaln #(12) e3176(.a(buffered_input), .b(12'b110001101000), .eq(weq3176));
    equaln #(12) e3177(.a(buffered_input), .b(12'b110001101001), .eq(weq3177));
    equaln #(12) e3178(.a(buffered_input), .b(12'b110001101010), .eq(weq3178));
    equaln #(12) e3179(.a(buffered_input), .b(12'b110001101011), .eq(weq3179));
    equaln #(12) e3180(.a(buffered_input), .b(12'b110001101100), .eq(weq3180));
    equaln #(12) e3181(.a(buffered_input), .b(12'b110001101101), .eq(weq3181));
    equaln #(12) e3182(.a(buffered_input), .b(12'b110001101110), .eq(weq3182));
    equaln #(12) e3183(.a(buffered_input), .b(12'b110001101111), .eq(weq3183));
    equaln #(12) e3184(.a(buffered_input), .b(12'b110001110000), .eq(weq3184));
    equaln #(12) e3185(.a(buffered_input), .b(12'b110001110001), .eq(weq3185));
    equaln #(12) e3186(.a(buffered_input), .b(12'b110001110010), .eq(weq3186));
    equaln #(12) e3187(.a(buffered_input), .b(12'b110001110011), .eq(weq3187));
    equaln #(12) e3188(.a(buffered_input), .b(12'b110001110100), .eq(weq3188));
    equaln #(12) e3189(.a(buffered_input), .b(12'b110001110101), .eq(weq3189));
    equaln #(12) e3190(.a(buffered_input), .b(12'b110001110110), .eq(weq3190));
    equaln #(12) e3191(.a(buffered_input), .b(12'b110001110111), .eq(weq3191));
    equaln #(12) e3192(.a(buffered_input), .b(12'b110001111000), .eq(weq3192));
    equaln #(12) e3193(.a(buffered_input), .b(12'b110001111001), .eq(weq3193));
    equaln #(12) e3194(.a(buffered_input), .b(12'b110001111010), .eq(weq3194));
    equaln #(12) e3195(.a(buffered_input), .b(12'b110001111011), .eq(weq3195));
    equaln #(12) e3196(.a(buffered_input), .b(12'b110001111100), .eq(weq3196));
    equaln #(12) e3197(.a(buffered_input), .b(12'b110001111101), .eq(weq3197));
    equaln #(12) e3198(.a(buffered_input), .b(12'b110001111110), .eq(weq3198));
    equaln #(12) e3199(.a(buffered_input), .b(12'b110001111111), .eq(weq3199));
    equaln #(12) e3200(.a(buffered_input), .b(12'b110010000000), .eq(weq3200));
    equaln #(12) e3201(.a(buffered_input), .b(12'b110010000001), .eq(weq3201));
    equaln #(12) e3202(.a(buffered_input), .b(12'b110010000010), .eq(weq3202));
    equaln #(12) e3203(.a(buffered_input), .b(12'b110010000011), .eq(weq3203));
    equaln #(12) e3204(.a(buffered_input), .b(12'b110010000100), .eq(weq3204));
    equaln #(12) e3205(.a(buffered_input), .b(12'b110010000101), .eq(weq3205));
    equaln #(12) e3206(.a(buffered_input), .b(12'b110010000110), .eq(weq3206));
    equaln #(12) e3207(.a(buffered_input), .b(12'b110010000111), .eq(weq3207));
    equaln #(12) e3208(.a(buffered_input), .b(12'b110010001000), .eq(weq3208));
    equaln #(12) e3209(.a(buffered_input), .b(12'b110010001001), .eq(weq3209));
    equaln #(12) e3210(.a(buffered_input), .b(12'b110010001010), .eq(weq3210));
    equaln #(12) e3211(.a(buffered_input), .b(12'b110010001011), .eq(weq3211));
    equaln #(12) e3212(.a(buffered_input), .b(12'b110010001100), .eq(weq3212));
    equaln #(12) e3213(.a(buffered_input), .b(12'b110010001101), .eq(weq3213));
    equaln #(12) e3214(.a(buffered_input), .b(12'b110010001110), .eq(weq3214));
    equaln #(12) e3215(.a(buffered_input), .b(12'b110010001111), .eq(weq3215));
    equaln #(12) e3216(.a(buffered_input), .b(12'b110010010000), .eq(weq3216));
    equaln #(12) e3217(.a(buffered_input), .b(12'b110010010001), .eq(weq3217));
    equaln #(12) e3218(.a(buffered_input), .b(12'b110010010010), .eq(weq3218));
    equaln #(12) e3219(.a(buffered_input), .b(12'b110010010011), .eq(weq3219));
    equaln #(12) e3220(.a(buffered_input), .b(12'b110010010100), .eq(weq3220));
    equaln #(12) e3221(.a(buffered_input), .b(12'b110010010101), .eq(weq3221));
    equaln #(12) e3222(.a(buffered_input), .b(12'b110010010110), .eq(weq3222));
    equaln #(12) e3223(.a(buffered_input), .b(12'b110010010111), .eq(weq3223));
    equaln #(12) e3224(.a(buffered_input), .b(12'b110010011000), .eq(weq3224));
    equaln #(12) e3225(.a(buffered_input), .b(12'b110010011001), .eq(weq3225));
    equaln #(12) e3226(.a(buffered_input), .b(12'b110010011010), .eq(weq3226));
    equaln #(12) e3227(.a(buffered_input), .b(12'b110010011011), .eq(weq3227));
    equaln #(12) e3228(.a(buffered_input), .b(12'b110010011100), .eq(weq3228));
    equaln #(12) e3229(.a(buffered_input), .b(12'b110010011101), .eq(weq3229));
    equaln #(12) e3230(.a(buffered_input), .b(12'b110010011110), .eq(weq3230));
    equaln #(12) e3231(.a(buffered_input), .b(12'b110010011111), .eq(weq3231));
    equaln #(12) e3232(.a(buffered_input), .b(12'b110010100000), .eq(weq3232));
    equaln #(12) e3233(.a(buffered_input), .b(12'b110010100001), .eq(weq3233));
    equaln #(12) e3234(.a(buffered_input), .b(12'b110010100010), .eq(weq3234));
    equaln #(12) e3235(.a(buffered_input), .b(12'b110010100011), .eq(weq3235));
    equaln #(12) e3236(.a(buffered_input), .b(12'b110010100100), .eq(weq3236));
    equaln #(12) e3237(.a(buffered_input), .b(12'b110010100101), .eq(weq3237));
    equaln #(12) e3238(.a(buffered_input), .b(12'b110010100110), .eq(weq3238));
    equaln #(12) e3239(.a(buffered_input), .b(12'b110010100111), .eq(weq3239));
    equaln #(12) e3240(.a(buffered_input), .b(12'b110010101000), .eq(weq3240));
    equaln #(12) e3241(.a(buffered_input), .b(12'b110010101001), .eq(weq3241));
    equaln #(12) e3242(.a(buffered_input), .b(12'b110010101010), .eq(weq3242));
    equaln #(12) e3243(.a(buffered_input), .b(12'b110010101011), .eq(weq3243));
    equaln #(12) e3244(.a(buffered_input), .b(12'b110010101100), .eq(weq3244));
    equaln #(12) e3245(.a(buffered_input), .b(12'b110010101101), .eq(weq3245));
    equaln #(12) e3246(.a(buffered_input), .b(12'b110010101110), .eq(weq3246));
    equaln #(12) e3247(.a(buffered_input), .b(12'b110010101111), .eq(weq3247));
    equaln #(12) e3248(.a(buffered_input), .b(12'b110010110000), .eq(weq3248));
    equaln #(12) e3249(.a(buffered_input), .b(12'b110010110001), .eq(weq3249));
    equaln #(12) e3250(.a(buffered_input), .b(12'b110010110010), .eq(weq3250));
    equaln #(12) e3251(.a(buffered_input), .b(12'b110010110011), .eq(weq3251));
    equaln #(12) e3252(.a(buffered_input), .b(12'b110010110100), .eq(weq3252));
    equaln #(12) e3253(.a(buffered_input), .b(12'b110010110101), .eq(weq3253));
    equaln #(12) e3254(.a(buffered_input), .b(12'b110010110110), .eq(weq3254));
    equaln #(12) e3255(.a(buffered_input), .b(12'b110010110111), .eq(weq3255));
    equaln #(12) e3256(.a(buffered_input), .b(12'b110010111000), .eq(weq3256));
    equaln #(12) e3257(.a(buffered_input), .b(12'b110010111001), .eq(weq3257));
    equaln #(12) e3258(.a(buffered_input), .b(12'b110010111010), .eq(weq3258));
    equaln #(12) e3259(.a(buffered_input), .b(12'b110010111011), .eq(weq3259));
    equaln #(12) e3260(.a(buffered_input), .b(12'b110010111100), .eq(weq3260));
    equaln #(12) e3261(.a(buffered_input), .b(12'b110010111101), .eq(weq3261));
    equaln #(12) e3262(.a(buffered_input), .b(12'b110010111110), .eq(weq3262));
    equaln #(12) e3263(.a(buffered_input), .b(12'b110010111111), .eq(weq3263));
    equaln #(12) e3264(.a(buffered_input), .b(12'b110011000000), .eq(weq3264));
    equaln #(12) e3265(.a(buffered_input), .b(12'b110011000001), .eq(weq3265));
    equaln #(12) e3266(.a(buffered_input), .b(12'b110011000010), .eq(weq3266));
    equaln #(12) e3267(.a(buffered_input), .b(12'b110011000011), .eq(weq3267));
    equaln #(12) e3268(.a(buffered_input), .b(12'b110011000100), .eq(weq3268));
    equaln #(12) e3269(.a(buffered_input), .b(12'b110011000101), .eq(weq3269));
    equaln #(12) e3270(.a(buffered_input), .b(12'b110011000110), .eq(weq3270));
    equaln #(12) e3271(.a(buffered_input), .b(12'b110011000111), .eq(weq3271));
    equaln #(12) e3272(.a(buffered_input), .b(12'b110011001000), .eq(weq3272));
    equaln #(12) e3273(.a(buffered_input), .b(12'b110011001001), .eq(weq3273));
    equaln #(12) e3274(.a(buffered_input), .b(12'b110011001010), .eq(weq3274));
    equaln #(12) e3275(.a(buffered_input), .b(12'b110011001011), .eq(weq3275));
    equaln #(12) e3276(.a(buffered_input), .b(12'b110011001100), .eq(weq3276));
    equaln #(12) e3277(.a(buffered_input), .b(12'b110011001101), .eq(weq3277));
    equaln #(12) e3278(.a(buffered_input), .b(12'b110011001110), .eq(weq3278));
    equaln #(12) e3279(.a(buffered_input), .b(12'b110011001111), .eq(weq3279));
    equaln #(12) e3280(.a(buffered_input), .b(12'b110011010000), .eq(weq3280));
    equaln #(12) e3281(.a(buffered_input), .b(12'b110011010001), .eq(weq3281));
    equaln #(12) e3282(.a(buffered_input), .b(12'b110011010010), .eq(weq3282));
    equaln #(12) e3283(.a(buffered_input), .b(12'b110011010011), .eq(weq3283));
    equaln #(12) e3284(.a(buffered_input), .b(12'b110011010100), .eq(weq3284));
    equaln #(12) e3285(.a(buffered_input), .b(12'b110011010101), .eq(weq3285));
    equaln #(12) e3286(.a(buffered_input), .b(12'b110011010110), .eq(weq3286));
    equaln #(12) e3287(.a(buffered_input), .b(12'b110011010111), .eq(weq3287));
    equaln #(12) e3288(.a(buffered_input), .b(12'b110011011000), .eq(weq3288));
    equaln #(12) e3289(.a(buffered_input), .b(12'b110011011001), .eq(weq3289));
    equaln #(12) e3290(.a(buffered_input), .b(12'b110011011010), .eq(weq3290));
    equaln #(12) e3291(.a(buffered_input), .b(12'b110011011011), .eq(weq3291));
    equaln #(12) e3292(.a(buffered_input), .b(12'b110011011100), .eq(weq3292));
    equaln #(12) e3293(.a(buffered_input), .b(12'b110011011101), .eq(weq3293));
    equaln #(12) e3294(.a(buffered_input), .b(12'b110011011110), .eq(weq3294));
    equaln #(12) e3295(.a(buffered_input), .b(12'b110011011111), .eq(weq3295));
    equaln #(12) e3296(.a(buffered_input), .b(12'b110011100000), .eq(weq3296));
    equaln #(12) e3297(.a(buffered_input), .b(12'b110011100001), .eq(weq3297));
    equaln #(12) e3298(.a(buffered_input), .b(12'b110011100010), .eq(weq3298));
    equaln #(12) e3299(.a(buffered_input), .b(12'b110011100011), .eq(weq3299));
    equaln #(12) e3300(.a(buffered_input), .b(12'b110011100100), .eq(weq3300));
    equaln #(12) e3301(.a(buffered_input), .b(12'b110011100101), .eq(weq3301));
    equaln #(12) e3302(.a(buffered_input), .b(12'b110011100110), .eq(weq3302));
    equaln #(12) e3303(.a(buffered_input), .b(12'b110011100111), .eq(weq3303));
    equaln #(12) e3304(.a(buffered_input), .b(12'b110011101000), .eq(weq3304));
    equaln #(12) e3305(.a(buffered_input), .b(12'b110011101001), .eq(weq3305));
    equaln #(12) e3306(.a(buffered_input), .b(12'b110011101010), .eq(weq3306));
    equaln #(12) e3307(.a(buffered_input), .b(12'b110011101011), .eq(weq3307));
    equaln #(12) e3308(.a(buffered_input), .b(12'b110011101100), .eq(weq3308));
    equaln #(12) e3309(.a(buffered_input), .b(12'b110011101101), .eq(weq3309));
    equaln #(12) e3310(.a(buffered_input), .b(12'b110011101110), .eq(weq3310));
    equaln #(12) e3311(.a(buffered_input), .b(12'b110011101111), .eq(weq3311));
    equaln #(12) e3312(.a(buffered_input), .b(12'b110011110000), .eq(weq3312));
    equaln #(12) e3313(.a(buffered_input), .b(12'b110011110001), .eq(weq3313));
    equaln #(12) e3314(.a(buffered_input), .b(12'b110011110010), .eq(weq3314));
    equaln #(12) e3315(.a(buffered_input), .b(12'b110011110011), .eq(weq3315));
    equaln #(12) e3316(.a(buffered_input), .b(12'b110011110100), .eq(weq3316));
    equaln #(12) e3317(.a(buffered_input), .b(12'b110011110101), .eq(weq3317));
    equaln #(12) e3318(.a(buffered_input), .b(12'b110011110110), .eq(weq3318));
    equaln #(12) e3319(.a(buffered_input), .b(12'b110011110111), .eq(weq3319));
    equaln #(12) e3320(.a(buffered_input), .b(12'b110011111000), .eq(weq3320));
    equaln #(12) e3321(.a(buffered_input), .b(12'b110011111001), .eq(weq3321));
    equaln #(12) e3322(.a(buffered_input), .b(12'b110011111010), .eq(weq3322));
    equaln #(12) e3323(.a(buffered_input), .b(12'b110011111011), .eq(weq3323));
    equaln #(12) e3324(.a(buffered_input), .b(12'b110011111100), .eq(weq3324));
    equaln #(12) e3325(.a(buffered_input), .b(12'b110011111101), .eq(weq3325));
    equaln #(12) e3326(.a(buffered_input), .b(12'b110011111110), .eq(weq3326));
    equaln #(12) e3327(.a(buffered_input), .b(12'b110011111111), .eq(weq3327));
    equaln #(12) e3328(.a(buffered_input), .b(12'b110100000000), .eq(weq3328));
    equaln #(12) e3329(.a(buffered_input), .b(12'b110100000001), .eq(weq3329));
    equaln #(12) e3330(.a(buffered_input), .b(12'b110100000010), .eq(weq3330));
    equaln #(12) e3331(.a(buffered_input), .b(12'b110100000011), .eq(weq3331));
    equaln #(12) e3332(.a(buffered_input), .b(12'b110100000100), .eq(weq3332));
    equaln #(12) e3333(.a(buffered_input), .b(12'b110100000101), .eq(weq3333));
    equaln #(12) e3334(.a(buffered_input), .b(12'b110100000110), .eq(weq3334));
    equaln #(12) e3335(.a(buffered_input), .b(12'b110100000111), .eq(weq3335));
    equaln #(12) e3336(.a(buffered_input), .b(12'b110100001000), .eq(weq3336));
    equaln #(12) e3337(.a(buffered_input), .b(12'b110100001001), .eq(weq3337));
    equaln #(12) e3338(.a(buffered_input), .b(12'b110100001010), .eq(weq3338));
    equaln #(12) e3339(.a(buffered_input), .b(12'b110100001011), .eq(weq3339));
    equaln #(12) e3340(.a(buffered_input), .b(12'b110100001100), .eq(weq3340));
    equaln #(12) e3341(.a(buffered_input), .b(12'b110100001101), .eq(weq3341));
    equaln #(12) e3342(.a(buffered_input), .b(12'b110100001110), .eq(weq3342));
    equaln #(12) e3343(.a(buffered_input), .b(12'b110100001111), .eq(weq3343));
    equaln #(12) e3344(.a(buffered_input), .b(12'b110100010000), .eq(weq3344));
    equaln #(12) e3345(.a(buffered_input), .b(12'b110100010001), .eq(weq3345));
    equaln #(12) e3346(.a(buffered_input), .b(12'b110100010010), .eq(weq3346));
    equaln #(12) e3347(.a(buffered_input), .b(12'b110100010011), .eq(weq3347));
    equaln #(12) e3348(.a(buffered_input), .b(12'b110100010100), .eq(weq3348));
    equaln #(12) e3349(.a(buffered_input), .b(12'b110100010101), .eq(weq3349));
    equaln #(12) e3350(.a(buffered_input), .b(12'b110100010110), .eq(weq3350));
    equaln #(12) e3351(.a(buffered_input), .b(12'b110100010111), .eq(weq3351));
    equaln #(12) e3352(.a(buffered_input), .b(12'b110100011000), .eq(weq3352));
    equaln #(12) e3353(.a(buffered_input), .b(12'b110100011001), .eq(weq3353));
    equaln #(12) e3354(.a(buffered_input), .b(12'b110100011010), .eq(weq3354));
    equaln #(12) e3355(.a(buffered_input), .b(12'b110100011011), .eq(weq3355));
    equaln #(12) e3356(.a(buffered_input), .b(12'b110100011100), .eq(weq3356));
    equaln #(12) e3357(.a(buffered_input), .b(12'b110100011101), .eq(weq3357));
    equaln #(12) e3358(.a(buffered_input), .b(12'b110100011110), .eq(weq3358));
    equaln #(12) e3359(.a(buffered_input), .b(12'b110100011111), .eq(weq3359));
    equaln #(12) e3360(.a(buffered_input), .b(12'b110100100000), .eq(weq3360));
    equaln #(12) e3361(.a(buffered_input), .b(12'b110100100001), .eq(weq3361));
    equaln #(12) e3362(.a(buffered_input), .b(12'b110100100010), .eq(weq3362));
    equaln #(12) e3363(.a(buffered_input), .b(12'b110100100011), .eq(weq3363));
    equaln #(12) e3364(.a(buffered_input), .b(12'b110100100100), .eq(weq3364));
    equaln #(12) e3365(.a(buffered_input), .b(12'b110100100101), .eq(weq3365));
    equaln #(12) e3366(.a(buffered_input), .b(12'b110100100110), .eq(weq3366));
    equaln #(12) e3367(.a(buffered_input), .b(12'b110100100111), .eq(weq3367));
    equaln #(12) e3368(.a(buffered_input), .b(12'b110100101000), .eq(weq3368));
    equaln #(12) e3369(.a(buffered_input), .b(12'b110100101001), .eq(weq3369));
    equaln #(12) e3370(.a(buffered_input), .b(12'b110100101010), .eq(weq3370));
    equaln #(12) e3371(.a(buffered_input), .b(12'b110100101011), .eq(weq3371));
    equaln #(12) e3372(.a(buffered_input), .b(12'b110100101100), .eq(weq3372));
    equaln #(12) e3373(.a(buffered_input), .b(12'b110100101101), .eq(weq3373));
    equaln #(12) e3374(.a(buffered_input), .b(12'b110100101110), .eq(weq3374));
    equaln #(12) e3375(.a(buffered_input), .b(12'b110100101111), .eq(weq3375));
    equaln #(12) e3376(.a(buffered_input), .b(12'b110100110000), .eq(weq3376));
    equaln #(12) e3377(.a(buffered_input), .b(12'b110100110001), .eq(weq3377));
    equaln #(12) e3378(.a(buffered_input), .b(12'b110100110010), .eq(weq3378));
    equaln #(12) e3379(.a(buffered_input), .b(12'b110100110011), .eq(weq3379));
    equaln #(12) e3380(.a(buffered_input), .b(12'b110100110100), .eq(weq3380));
    equaln #(12) e3381(.a(buffered_input), .b(12'b110100110101), .eq(weq3381));
    equaln #(12) e3382(.a(buffered_input), .b(12'b110100110110), .eq(weq3382));
    equaln #(12) e3383(.a(buffered_input), .b(12'b110100110111), .eq(weq3383));
    equaln #(12) e3384(.a(buffered_input), .b(12'b110100111000), .eq(weq3384));
    equaln #(12) e3385(.a(buffered_input), .b(12'b110100111001), .eq(weq3385));
    equaln #(12) e3386(.a(buffered_input), .b(12'b110100111010), .eq(weq3386));
    equaln #(12) e3387(.a(buffered_input), .b(12'b110100111011), .eq(weq3387));
    equaln #(12) e3388(.a(buffered_input), .b(12'b110100111100), .eq(weq3388));
    equaln #(12) e3389(.a(buffered_input), .b(12'b110100111101), .eq(weq3389));
    equaln #(12) e3390(.a(buffered_input), .b(12'b110100111110), .eq(weq3390));
    equaln #(12) e3391(.a(buffered_input), .b(12'b110100111111), .eq(weq3391));
    equaln #(12) e3392(.a(buffered_input), .b(12'b110101000000), .eq(weq3392));
    equaln #(12) e3393(.a(buffered_input), .b(12'b110101000001), .eq(weq3393));
    equaln #(12) e3394(.a(buffered_input), .b(12'b110101000010), .eq(weq3394));
    equaln #(12) e3395(.a(buffered_input), .b(12'b110101000011), .eq(weq3395));
    equaln #(12) e3396(.a(buffered_input), .b(12'b110101000100), .eq(weq3396));
    equaln #(12) e3397(.a(buffered_input), .b(12'b110101000101), .eq(weq3397));
    equaln #(12) e3398(.a(buffered_input), .b(12'b110101000110), .eq(weq3398));
    equaln #(12) e3399(.a(buffered_input), .b(12'b110101000111), .eq(weq3399));
    equaln #(12) e3400(.a(buffered_input), .b(12'b110101001000), .eq(weq3400));
    equaln #(12) e3401(.a(buffered_input), .b(12'b110101001001), .eq(weq3401));
    equaln #(12) e3402(.a(buffered_input), .b(12'b110101001010), .eq(weq3402));
    equaln #(12) e3403(.a(buffered_input), .b(12'b110101001011), .eq(weq3403));
    equaln #(12) e3404(.a(buffered_input), .b(12'b110101001100), .eq(weq3404));
    equaln #(12) e3405(.a(buffered_input), .b(12'b110101001101), .eq(weq3405));
    equaln #(12) e3406(.a(buffered_input), .b(12'b110101001110), .eq(weq3406));
    equaln #(12) e3407(.a(buffered_input), .b(12'b110101001111), .eq(weq3407));
    equaln #(12) e3408(.a(buffered_input), .b(12'b110101010000), .eq(weq3408));
    equaln #(12) e3409(.a(buffered_input), .b(12'b110101010001), .eq(weq3409));
    equaln #(12) e3410(.a(buffered_input), .b(12'b110101010010), .eq(weq3410));
    equaln #(12) e3411(.a(buffered_input), .b(12'b110101010011), .eq(weq3411));
    equaln #(12) e3412(.a(buffered_input), .b(12'b110101010100), .eq(weq3412));
    equaln #(12) e3413(.a(buffered_input), .b(12'b110101010101), .eq(weq3413));
    equaln #(12) e3414(.a(buffered_input), .b(12'b110101010110), .eq(weq3414));
    equaln #(12) e3415(.a(buffered_input), .b(12'b110101010111), .eq(weq3415));
    equaln #(12) e3416(.a(buffered_input), .b(12'b110101011000), .eq(weq3416));
    equaln #(12) e3417(.a(buffered_input), .b(12'b110101011001), .eq(weq3417));
    equaln #(12) e3418(.a(buffered_input), .b(12'b110101011010), .eq(weq3418));
    equaln #(12) e3419(.a(buffered_input), .b(12'b110101011011), .eq(weq3419));
    equaln #(12) e3420(.a(buffered_input), .b(12'b110101011100), .eq(weq3420));
    equaln #(12) e3421(.a(buffered_input), .b(12'b110101011101), .eq(weq3421));
    equaln #(12) e3422(.a(buffered_input), .b(12'b110101011110), .eq(weq3422));
    equaln #(12) e3423(.a(buffered_input), .b(12'b110101011111), .eq(weq3423));
    equaln #(12) e3424(.a(buffered_input), .b(12'b110101100000), .eq(weq3424));
    equaln #(12) e3425(.a(buffered_input), .b(12'b110101100001), .eq(weq3425));
    equaln #(12) e3426(.a(buffered_input), .b(12'b110101100010), .eq(weq3426));
    equaln #(12) e3427(.a(buffered_input), .b(12'b110101100011), .eq(weq3427));
    equaln #(12) e3428(.a(buffered_input), .b(12'b110101100100), .eq(weq3428));
    equaln #(12) e3429(.a(buffered_input), .b(12'b110101100101), .eq(weq3429));
    equaln #(12) e3430(.a(buffered_input), .b(12'b110101100110), .eq(weq3430));
    equaln #(12) e3431(.a(buffered_input), .b(12'b110101100111), .eq(weq3431));
    equaln #(12) e3432(.a(buffered_input), .b(12'b110101101000), .eq(weq3432));
    equaln #(12) e3433(.a(buffered_input), .b(12'b110101101001), .eq(weq3433));
    equaln #(12) e3434(.a(buffered_input), .b(12'b110101101010), .eq(weq3434));
    equaln #(12) e3435(.a(buffered_input), .b(12'b110101101011), .eq(weq3435));
    equaln #(12) e3436(.a(buffered_input), .b(12'b110101101100), .eq(weq3436));
    equaln #(12) e3437(.a(buffered_input), .b(12'b110101101101), .eq(weq3437));
    equaln #(12) e3438(.a(buffered_input), .b(12'b110101101110), .eq(weq3438));
    equaln #(12) e3439(.a(buffered_input), .b(12'b110101101111), .eq(weq3439));
    equaln #(12) e3440(.a(buffered_input), .b(12'b110101110000), .eq(weq3440));
    equaln #(12) e3441(.a(buffered_input), .b(12'b110101110001), .eq(weq3441));
    equaln #(12) e3442(.a(buffered_input), .b(12'b110101110010), .eq(weq3442));
    equaln #(12) e3443(.a(buffered_input), .b(12'b110101110011), .eq(weq3443));
    equaln #(12) e3444(.a(buffered_input), .b(12'b110101110100), .eq(weq3444));
    equaln #(12) e3445(.a(buffered_input), .b(12'b110101110101), .eq(weq3445));
    equaln #(12) e3446(.a(buffered_input), .b(12'b110101110110), .eq(weq3446));
    equaln #(12) e3447(.a(buffered_input), .b(12'b110101110111), .eq(weq3447));
    equaln #(12) e3448(.a(buffered_input), .b(12'b110101111000), .eq(weq3448));
    equaln #(12) e3449(.a(buffered_input), .b(12'b110101111001), .eq(weq3449));
    equaln #(12) e3450(.a(buffered_input), .b(12'b110101111010), .eq(weq3450));
    equaln #(12) e3451(.a(buffered_input), .b(12'b110101111011), .eq(weq3451));
    equaln #(12) e3452(.a(buffered_input), .b(12'b110101111100), .eq(weq3452));
    equaln #(12) e3453(.a(buffered_input), .b(12'b110101111101), .eq(weq3453));
    equaln #(12) e3454(.a(buffered_input), .b(12'b110101111110), .eq(weq3454));
    equaln #(12) e3455(.a(buffered_input), .b(12'b110101111111), .eq(weq3455));
    equaln #(12) e3456(.a(buffered_input), .b(12'b110110000000), .eq(weq3456));
    equaln #(12) e3457(.a(buffered_input), .b(12'b110110000001), .eq(weq3457));
    equaln #(12) e3458(.a(buffered_input), .b(12'b110110000010), .eq(weq3458));
    equaln #(12) e3459(.a(buffered_input), .b(12'b110110000011), .eq(weq3459));
    equaln #(12) e3460(.a(buffered_input), .b(12'b110110000100), .eq(weq3460));
    equaln #(12) e3461(.a(buffered_input), .b(12'b110110000101), .eq(weq3461));
    equaln #(12) e3462(.a(buffered_input), .b(12'b110110000110), .eq(weq3462));
    equaln #(12) e3463(.a(buffered_input), .b(12'b110110000111), .eq(weq3463));
    equaln #(12) e3464(.a(buffered_input), .b(12'b110110001000), .eq(weq3464));
    equaln #(12) e3465(.a(buffered_input), .b(12'b110110001001), .eq(weq3465));
    equaln #(12) e3466(.a(buffered_input), .b(12'b110110001010), .eq(weq3466));
    equaln #(12) e3467(.a(buffered_input), .b(12'b110110001011), .eq(weq3467));
    equaln #(12) e3468(.a(buffered_input), .b(12'b110110001100), .eq(weq3468));
    equaln #(12) e3469(.a(buffered_input), .b(12'b110110001101), .eq(weq3469));
    equaln #(12) e3470(.a(buffered_input), .b(12'b110110001110), .eq(weq3470));
    equaln #(12) e3471(.a(buffered_input), .b(12'b110110001111), .eq(weq3471));
    equaln #(12) e3472(.a(buffered_input), .b(12'b110110010000), .eq(weq3472));
    equaln #(12) e3473(.a(buffered_input), .b(12'b110110010001), .eq(weq3473));
    equaln #(12) e3474(.a(buffered_input), .b(12'b110110010010), .eq(weq3474));
    equaln #(12) e3475(.a(buffered_input), .b(12'b110110010011), .eq(weq3475));
    equaln #(12) e3476(.a(buffered_input), .b(12'b110110010100), .eq(weq3476));
    equaln #(12) e3477(.a(buffered_input), .b(12'b110110010101), .eq(weq3477));
    equaln #(12) e3478(.a(buffered_input), .b(12'b110110010110), .eq(weq3478));
    equaln #(12) e3479(.a(buffered_input), .b(12'b110110010111), .eq(weq3479));
    equaln #(12) e3480(.a(buffered_input), .b(12'b110110011000), .eq(weq3480));
    equaln #(12) e3481(.a(buffered_input), .b(12'b110110011001), .eq(weq3481));
    equaln #(12) e3482(.a(buffered_input), .b(12'b110110011010), .eq(weq3482));
    equaln #(12) e3483(.a(buffered_input), .b(12'b110110011011), .eq(weq3483));
    equaln #(12) e3484(.a(buffered_input), .b(12'b110110011100), .eq(weq3484));
    equaln #(12) e3485(.a(buffered_input), .b(12'b110110011101), .eq(weq3485));
    equaln #(12) e3486(.a(buffered_input), .b(12'b110110011110), .eq(weq3486));
    equaln #(12) e3487(.a(buffered_input), .b(12'b110110011111), .eq(weq3487));
    equaln #(12) e3488(.a(buffered_input), .b(12'b110110100000), .eq(weq3488));
    equaln #(12) e3489(.a(buffered_input), .b(12'b110110100001), .eq(weq3489));
    equaln #(12) e3490(.a(buffered_input), .b(12'b110110100010), .eq(weq3490));
    equaln #(12) e3491(.a(buffered_input), .b(12'b110110100011), .eq(weq3491));
    equaln #(12) e3492(.a(buffered_input), .b(12'b110110100100), .eq(weq3492));
    equaln #(12) e3493(.a(buffered_input), .b(12'b110110100101), .eq(weq3493));
    equaln #(12) e3494(.a(buffered_input), .b(12'b110110100110), .eq(weq3494));
    equaln #(12) e3495(.a(buffered_input), .b(12'b110110100111), .eq(weq3495));
    equaln #(12) e3496(.a(buffered_input), .b(12'b110110101000), .eq(weq3496));
    equaln #(12) e3497(.a(buffered_input), .b(12'b110110101001), .eq(weq3497));
    equaln #(12) e3498(.a(buffered_input), .b(12'b110110101010), .eq(weq3498));
    equaln #(12) e3499(.a(buffered_input), .b(12'b110110101011), .eq(weq3499));
    equaln #(12) e3500(.a(buffered_input), .b(12'b110110101100), .eq(weq3500));
    equaln #(12) e3501(.a(buffered_input), .b(12'b110110101101), .eq(weq3501));
    equaln #(12) e3502(.a(buffered_input), .b(12'b110110101110), .eq(weq3502));
    equaln #(12) e3503(.a(buffered_input), .b(12'b110110101111), .eq(weq3503));
    equaln #(12) e3504(.a(buffered_input), .b(12'b110110110000), .eq(weq3504));
    equaln #(12) e3505(.a(buffered_input), .b(12'b110110110001), .eq(weq3505));
    equaln #(12) e3506(.a(buffered_input), .b(12'b110110110010), .eq(weq3506));
    equaln #(12) e3507(.a(buffered_input), .b(12'b110110110011), .eq(weq3507));
    equaln #(12) e3508(.a(buffered_input), .b(12'b110110110100), .eq(weq3508));
    equaln #(12) e3509(.a(buffered_input), .b(12'b110110110101), .eq(weq3509));
    equaln #(12) e3510(.a(buffered_input), .b(12'b110110110110), .eq(weq3510));
    equaln #(12) e3511(.a(buffered_input), .b(12'b110110110111), .eq(weq3511));
    equaln #(12) e3512(.a(buffered_input), .b(12'b110110111000), .eq(weq3512));
    equaln #(12) e3513(.a(buffered_input), .b(12'b110110111001), .eq(weq3513));
    equaln #(12) e3514(.a(buffered_input), .b(12'b110110111010), .eq(weq3514));
    equaln #(12) e3515(.a(buffered_input), .b(12'b110110111011), .eq(weq3515));
    equaln #(12) e3516(.a(buffered_input), .b(12'b110110111100), .eq(weq3516));
    equaln #(12) e3517(.a(buffered_input), .b(12'b110110111101), .eq(weq3517));
    equaln #(12) e3518(.a(buffered_input), .b(12'b110110111110), .eq(weq3518));
    equaln #(12) e3519(.a(buffered_input), .b(12'b110110111111), .eq(weq3519));
    equaln #(12) e3520(.a(buffered_input), .b(12'b110111000000), .eq(weq3520));
    equaln #(12) e3521(.a(buffered_input), .b(12'b110111000001), .eq(weq3521));
    equaln #(12) e3522(.a(buffered_input), .b(12'b110111000010), .eq(weq3522));
    equaln #(12) e3523(.a(buffered_input), .b(12'b110111000011), .eq(weq3523));
    equaln #(12) e3524(.a(buffered_input), .b(12'b110111000100), .eq(weq3524));
    equaln #(12) e3525(.a(buffered_input), .b(12'b110111000101), .eq(weq3525));
    equaln #(12) e3526(.a(buffered_input), .b(12'b110111000110), .eq(weq3526));
    equaln #(12) e3527(.a(buffered_input), .b(12'b110111000111), .eq(weq3527));
    equaln #(12) e3528(.a(buffered_input), .b(12'b110111001000), .eq(weq3528));
    equaln #(12) e3529(.a(buffered_input), .b(12'b110111001001), .eq(weq3529));
    equaln #(12) e3530(.a(buffered_input), .b(12'b110111001010), .eq(weq3530));
    equaln #(12) e3531(.a(buffered_input), .b(12'b110111001011), .eq(weq3531));
    equaln #(12) e3532(.a(buffered_input), .b(12'b110111001100), .eq(weq3532));
    equaln #(12) e3533(.a(buffered_input), .b(12'b110111001101), .eq(weq3533));
    equaln #(12) e3534(.a(buffered_input), .b(12'b110111001110), .eq(weq3534));
    equaln #(12) e3535(.a(buffered_input), .b(12'b110111001111), .eq(weq3535));
    equaln #(12) e3536(.a(buffered_input), .b(12'b110111010000), .eq(weq3536));
    equaln #(12) e3537(.a(buffered_input), .b(12'b110111010001), .eq(weq3537));
    equaln #(12) e3538(.a(buffered_input), .b(12'b110111010010), .eq(weq3538));
    equaln #(12) e3539(.a(buffered_input), .b(12'b110111010011), .eq(weq3539));
    equaln #(12) e3540(.a(buffered_input), .b(12'b110111010100), .eq(weq3540));
    equaln #(12) e3541(.a(buffered_input), .b(12'b110111010101), .eq(weq3541));
    equaln #(12) e3542(.a(buffered_input), .b(12'b110111010110), .eq(weq3542));
    equaln #(12) e3543(.a(buffered_input), .b(12'b110111010111), .eq(weq3543));
    equaln #(12) e3544(.a(buffered_input), .b(12'b110111011000), .eq(weq3544));
    equaln #(12) e3545(.a(buffered_input), .b(12'b110111011001), .eq(weq3545));
    equaln #(12) e3546(.a(buffered_input), .b(12'b110111011010), .eq(weq3546));
    equaln #(12) e3547(.a(buffered_input), .b(12'b110111011011), .eq(weq3547));
    equaln #(12) e3548(.a(buffered_input), .b(12'b110111011100), .eq(weq3548));
    equaln #(12) e3549(.a(buffered_input), .b(12'b110111011101), .eq(weq3549));
    equaln #(12) e3550(.a(buffered_input), .b(12'b110111011110), .eq(weq3550));
    equaln #(12) e3551(.a(buffered_input), .b(12'b110111011111), .eq(weq3551));
    equaln #(12) e3552(.a(buffered_input), .b(12'b110111100000), .eq(weq3552));
    equaln #(12) e3553(.a(buffered_input), .b(12'b110111100001), .eq(weq3553));
    equaln #(12) e3554(.a(buffered_input), .b(12'b110111100010), .eq(weq3554));
    equaln #(12) e3555(.a(buffered_input), .b(12'b110111100011), .eq(weq3555));
    equaln #(12) e3556(.a(buffered_input), .b(12'b110111100100), .eq(weq3556));
    equaln #(12) e3557(.a(buffered_input), .b(12'b110111100101), .eq(weq3557));
    equaln #(12) e3558(.a(buffered_input), .b(12'b110111100110), .eq(weq3558));
    equaln #(12) e3559(.a(buffered_input), .b(12'b110111100111), .eq(weq3559));
    equaln #(12) e3560(.a(buffered_input), .b(12'b110111101000), .eq(weq3560));
    equaln #(12) e3561(.a(buffered_input), .b(12'b110111101001), .eq(weq3561));
    equaln #(12) e3562(.a(buffered_input), .b(12'b110111101010), .eq(weq3562));
    equaln #(12) e3563(.a(buffered_input), .b(12'b110111101011), .eq(weq3563));
    equaln #(12) e3564(.a(buffered_input), .b(12'b110111101100), .eq(weq3564));
    equaln #(12) e3565(.a(buffered_input), .b(12'b110111101101), .eq(weq3565));
    equaln #(12) e3566(.a(buffered_input), .b(12'b110111101110), .eq(weq3566));
    equaln #(12) e3567(.a(buffered_input), .b(12'b110111101111), .eq(weq3567));
    equaln #(12) e3568(.a(buffered_input), .b(12'b110111110000), .eq(weq3568));
    equaln #(12) e3569(.a(buffered_input), .b(12'b110111110001), .eq(weq3569));
    equaln #(12) e3570(.a(buffered_input), .b(12'b110111110010), .eq(weq3570));
    equaln #(12) e3571(.a(buffered_input), .b(12'b110111110011), .eq(weq3571));
    equaln #(12) e3572(.a(buffered_input), .b(12'b110111110100), .eq(weq3572));
    equaln #(12) e3573(.a(buffered_input), .b(12'b110111110101), .eq(weq3573));
    equaln #(12) e3574(.a(buffered_input), .b(12'b110111110110), .eq(weq3574));
    equaln #(12) e3575(.a(buffered_input), .b(12'b110111110111), .eq(weq3575));
    equaln #(12) e3576(.a(buffered_input), .b(12'b110111111000), .eq(weq3576));
    equaln #(12) e3577(.a(buffered_input), .b(12'b110111111001), .eq(weq3577));
    equaln #(12) e3578(.a(buffered_input), .b(12'b110111111010), .eq(weq3578));
    equaln #(12) e3579(.a(buffered_input), .b(12'b110111111011), .eq(weq3579));
    equaln #(12) e3580(.a(buffered_input), .b(12'b110111111100), .eq(weq3580));
    equaln #(12) e3581(.a(buffered_input), .b(12'b110111111101), .eq(weq3581));
    equaln #(12) e3582(.a(buffered_input), .b(12'b110111111110), .eq(weq3582));
    equaln #(12) e3583(.a(buffered_input), .b(12'b110111111111), .eq(weq3583));
    equaln #(12) e3584(.a(buffered_input), .b(12'b111000000000), .eq(weq3584));
    equaln #(12) e3585(.a(buffered_input), .b(12'b111000000001), .eq(weq3585));
    equaln #(12) e3586(.a(buffered_input), .b(12'b111000000010), .eq(weq3586));
    equaln #(12) e3587(.a(buffered_input), .b(12'b111000000011), .eq(weq3587));
    equaln #(12) e3588(.a(buffered_input), .b(12'b111000000100), .eq(weq3588));
    equaln #(12) e3589(.a(buffered_input), .b(12'b111000000101), .eq(weq3589));
    equaln #(12) e3590(.a(buffered_input), .b(12'b111000000110), .eq(weq3590));
    equaln #(12) e3591(.a(buffered_input), .b(12'b111000000111), .eq(weq3591));
    equaln #(12) e3592(.a(buffered_input), .b(12'b111000001000), .eq(weq3592));
    equaln #(12) e3593(.a(buffered_input), .b(12'b111000001001), .eq(weq3593));
    equaln #(12) e3594(.a(buffered_input), .b(12'b111000001010), .eq(weq3594));
    equaln #(12) e3595(.a(buffered_input), .b(12'b111000001011), .eq(weq3595));
    equaln #(12) e3596(.a(buffered_input), .b(12'b111000001100), .eq(weq3596));
    equaln #(12) e3597(.a(buffered_input), .b(12'b111000001101), .eq(weq3597));
    equaln #(12) e3598(.a(buffered_input), .b(12'b111000001110), .eq(weq3598));
    equaln #(12) e3599(.a(buffered_input), .b(12'b111000001111), .eq(weq3599));
    equaln #(12) e3600(.a(buffered_input), .b(12'b111000010000), .eq(weq3600));
    equaln #(12) e3601(.a(buffered_input), .b(12'b111000010001), .eq(weq3601));
    equaln #(12) e3602(.a(buffered_input), .b(12'b111000010010), .eq(weq3602));
    equaln #(12) e3603(.a(buffered_input), .b(12'b111000010011), .eq(weq3603));
    equaln #(12) e3604(.a(buffered_input), .b(12'b111000010100), .eq(weq3604));
    equaln #(12) e3605(.a(buffered_input), .b(12'b111000010101), .eq(weq3605));
    equaln #(12) e3606(.a(buffered_input), .b(12'b111000010110), .eq(weq3606));
    equaln #(12) e3607(.a(buffered_input), .b(12'b111000010111), .eq(weq3607));
    equaln #(12) e3608(.a(buffered_input), .b(12'b111000011000), .eq(weq3608));
    equaln #(12) e3609(.a(buffered_input), .b(12'b111000011001), .eq(weq3609));
    equaln #(12) e3610(.a(buffered_input), .b(12'b111000011010), .eq(weq3610));
    equaln #(12) e3611(.a(buffered_input), .b(12'b111000011011), .eq(weq3611));
    equaln #(12) e3612(.a(buffered_input), .b(12'b111000011100), .eq(weq3612));
    equaln #(12) e3613(.a(buffered_input), .b(12'b111000011101), .eq(weq3613));
    equaln #(12) e3614(.a(buffered_input), .b(12'b111000011110), .eq(weq3614));
    equaln #(12) e3615(.a(buffered_input), .b(12'b111000011111), .eq(weq3615));
    equaln #(12) e3616(.a(buffered_input), .b(12'b111000100000), .eq(weq3616));
    equaln #(12) e3617(.a(buffered_input), .b(12'b111000100001), .eq(weq3617));
    equaln #(12) e3618(.a(buffered_input), .b(12'b111000100010), .eq(weq3618));
    equaln #(12) e3619(.a(buffered_input), .b(12'b111000100011), .eq(weq3619));
    equaln #(12) e3620(.a(buffered_input), .b(12'b111000100100), .eq(weq3620));
    equaln #(12) e3621(.a(buffered_input), .b(12'b111000100101), .eq(weq3621));
    equaln #(12) e3622(.a(buffered_input), .b(12'b111000100110), .eq(weq3622));
    equaln #(12) e3623(.a(buffered_input), .b(12'b111000100111), .eq(weq3623));
    equaln #(12) e3624(.a(buffered_input), .b(12'b111000101000), .eq(weq3624));
    equaln #(12) e3625(.a(buffered_input), .b(12'b111000101001), .eq(weq3625));
    equaln #(12) e3626(.a(buffered_input), .b(12'b111000101010), .eq(weq3626));
    equaln #(12) e3627(.a(buffered_input), .b(12'b111000101011), .eq(weq3627));
    equaln #(12) e3628(.a(buffered_input), .b(12'b111000101100), .eq(weq3628));
    equaln #(12) e3629(.a(buffered_input), .b(12'b111000101101), .eq(weq3629));
    equaln #(12) e3630(.a(buffered_input), .b(12'b111000101110), .eq(weq3630));
    equaln #(12) e3631(.a(buffered_input), .b(12'b111000101111), .eq(weq3631));
    equaln #(12) e3632(.a(buffered_input), .b(12'b111000110000), .eq(weq3632));
    equaln #(12) e3633(.a(buffered_input), .b(12'b111000110001), .eq(weq3633));
    equaln #(12) e3634(.a(buffered_input), .b(12'b111000110010), .eq(weq3634));
    equaln #(12) e3635(.a(buffered_input), .b(12'b111000110011), .eq(weq3635));
    equaln #(12) e3636(.a(buffered_input), .b(12'b111000110100), .eq(weq3636));
    equaln #(12) e3637(.a(buffered_input), .b(12'b111000110101), .eq(weq3637));
    equaln #(12) e3638(.a(buffered_input), .b(12'b111000110110), .eq(weq3638));
    equaln #(12) e3639(.a(buffered_input), .b(12'b111000110111), .eq(weq3639));
    equaln #(12) e3640(.a(buffered_input), .b(12'b111000111000), .eq(weq3640));
    equaln #(12) e3641(.a(buffered_input), .b(12'b111000111001), .eq(weq3641));
    equaln #(12) e3642(.a(buffered_input), .b(12'b111000111010), .eq(weq3642));
    equaln #(12) e3643(.a(buffered_input), .b(12'b111000111011), .eq(weq3643));
    equaln #(12) e3644(.a(buffered_input), .b(12'b111000111100), .eq(weq3644));
    equaln #(12) e3645(.a(buffered_input), .b(12'b111000111101), .eq(weq3645));
    equaln #(12) e3646(.a(buffered_input), .b(12'b111000111110), .eq(weq3646));
    equaln #(12) e3647(.a(buffered_input), .b(12'b111000111111), .eq(weq3647));
    equaln #(12) e3648(.a(buffered_input), .b(12'b111001000000), .eq(weq3648));
    equaln #(12) e3649(.a(buffered_input), .b(12'b111001000001), .eq(weq3649));
    equaln #(12) e3650(.a(buffered_input), .b(12'b111001000010), .eq(weq3650));
    equaln #(12) e3651(.a(buffered_input), .b(12'b111001000011), .eq(weq3651));
    equaln #(12) e3652(.a(buffered_input), .b(12'b111001000100), .eq(weq3652));
    equaln #(12) e3653(.a(buffered_input), .b(12'b111001000101), .eq(weq3653));
    equaln #(12) e3654(.a(buffered_input), .b(12'b111001000110), .eq(weq3654));
    equaln #(12) e3655(.a(buffered_input), .b(12'b111001000111), .eq(weq3655));
    equaln #(12) e3656(.a(buffered_input), .b(12'b111001001000), .eq(weq3656));
    equaln #(12) e3657(.a(buffered_input), .b(12'b111001001001), .eq(weq3657));
    equaln #(12) e3658(.a(buffered_input), .b(12'b111001001010), .eq(weq3658));
    equaln #(12) e3659(.a(buffered_input), .b(12'b111001001011), .eq(weq3659));
    equaln #(12) e3660(.a(buffered_input), .b(12'b111001001100), .eq(weq3660));
    equaln #(12) e3661(.a(buffered_input), .b(12'b111001001101), .eq(weq3661));
    equaln #(12) e3662(.a(buffered_input), .b(12'b111001001110), .eq(weq3662));
    equaln #(12) e3663(.a(buffered_input), .b(12'b111001001111), .eq(weq3663));
    equaln #(12) e3664(.a(buffered_input), .b(12'b111001010000), .eq(weq3664));
    equaln #(12) e3665(.a(buffered_input), .b(12'b111001010001), .eq(weq3665));
    equaln #(12) e3666(.a(buffered_input), .b(12'b111001010010), .eq(weq3666));
    equaln #(12) e3667(.a(buffered_input), .b(12'b111001010011), .eq(weq3667));
    equaln #(12) e3668(.a(buffered_input), .b(12'b111001010100), .eq(weq3668));
    equaln #(12) e3669(.a(buffered_input), .b(12'b111001010101), .eq(weq3669));
    equaln #(12) e3670(.a(buffered_input), .b(12'b111001010110), .eq(weq3670));
    equaln #(12) e3671(.a(buffered_input), .b(12'b111001010111), .eq(weq3671));
    equaln #(12) e3672(.a(buffered_input), .b(12'b111001011000), .eq(weq3672));
    equaln #(12) e3673(.a(buffered_input), .b(12'b111001011001), .eq(weq3673));
    equaln #(12) e3674(.a(buffered_input), .b(12'b111001011010), .eq(weq3674));
    equaln #(12) e3675(.a(buffered_input), .b(12'b111001011011), .eq(weq3675));
    equaln #(12) e3676(.a(buffered_input), .b(12'b111001011100), .eq(weq3676));
    equaln #(12) e3677(.a(buffered_input), .b(12'b111001011101), .eq(weq3677));
    equaln #(12) e3678(.a(buffered_input), .b(12'b111001011110), .eq(weq3678));
    equaln #(12) e3679(.a(buffered_input), .b(12'b111001011111), .eq(weq3679));
    equaln #(12) e3680(.a(buffered_input), .b(12'b111001100000), .eq(weq3680));
    equaln #(12) e3681(.a(buffered_input), .b(12'b111001100001), .eq(weq3681));
    equaln #(12) e3682(.a(buffered_input), .b(12'b111001100010), .eq(weq3682));
    equaln #(12) e3683(.a(buffered_input), .b(12'b111001100011), .eq(weq3683));
    equaln #(12) e3684(.a(buffered_input), .b(12'b111001100100), .eq(weq3684));
    equaln #(12) e3685(.a(buffered_input), .b(12'b111001100101), .eq(weq3685));
    equaln #(12) e3686(.a(buffered_input), .b(12'b111001100110), .eq(weq3686));
    equaln #(12) e3687(.a(buffered_input), .b(12'b111001100111), .eq(weq3687));
    equaln #(12) e3688(.a(buffered_input), .b(12'b111001101000), .eq(weq3688));
    equaln #(12) e3689(.a(buffered_input), .b(12'b111001101001), .eq(weq3689));
    equaln #(12) e3690(.a(buffered_input), .b(12'b111001101010), .eq(weq3690));
    equaln #(12) e3691(.a(buffered_input), .b(12'b111001101011), .eq(weq3691));
    equaln #(12) e3692(.a(buffered_input), .b(12'b111001101100), .eq(weq3692));
    equaln #(12) e3693(.a(buffered_input), .b(12'b111001101101), .eq(weq3693));
    equaln #(12) e3694(.a(buffered_input), .b(12'b111001101110), .eq(weq3694));
    equaln #(12) e3695(.a(buffered_input), .b(12'b111001101111), .eq(weq3695));
    equaln #(12) e3696(.a(buffered_input), .b(12'b111001110000), .eq(weq3696));
    equaln #(12) e3697(.a(buffered_input), .b(12'b111001110001), .eq(weq3697));
    equaln #(12) e3698(.a(buffered_input), .b(12'b111001110010), .eq(weq3698));
    equaln #(12) e3699(.a(buffered_input), .b(12'b111001110011), .eq(weq3699));
    equaln #(12) e3700(.a(buffered_input), .b(12'b111001110100), .eq(weq3700));
    equaln #(12) e3701(.a(buffered_input), .b(12'b111001110101), .eq(weq3701));
    equaln #(12) e3702(.a(buffered_input), .b(12'b111001110110), .eq(weq3702));
    equaln #(12) e3703(.a(buffered_input), .b(12'b111001110111), .eq(weq3703));
    equaln #(12) e3704(.a(buffered_input), .b(12'b111001111000), .eq(weq3704));
    equaln #(12) e3705(.a(buffered_input), .b(12'b111001111001), .eq(weq3705));
    equaln #(12) e3706(.a(buffered_input), .b(12'b111001111010), .eq(weq3706));
    equaln #(12) e3707(.a(buffered_input), .b(12'b111001111011), .eq(weq3707));
    equaln #(12) e3708(.a(buffered_input), .b(12'b111001111100), .eq(weq3708));
    equaln #(12) e3709(.a(buffered_input), .b(12'b111001111101), .eq(weq3709));
    equaln #(12) e3710(.a(buffered_input), .b(12'b111001111110), .eq(weq3710));
    equaln #(12) e3711(.a(buffered_input), .b(12'b111001111111), .eq(weq3711));
    equaln #(12) e3712(.a(buffered_input), .b(12'b111010000000), .eq(weq3712));
    equaln #(12) e3713(.a(buffered_input), .b(12'b111010000001), .eq(weq3713));
    equaln #(12) e3714(.a(buffered_input), .b(12'b111010000010), .eq(weq3714));
    equaln #(12) e3715(.a(buffered_input), .b(12'b111010000011), .eq(weq3715));
    equaln #(12) e3716(.a(buffered_input), .b(12'b111010000100), .eq(weq3716));
    equaln #(12) e3717(.a(buffered_input), .b(12'b111010000101), .eq(weq3717));
    equaln #(12) e3718(.a(buffered_input), .b(12'b111010000110), .eq(weq3718));
    equaln #(12) e3719(.a(buffered_input), .b(12'b111010000111), .eq(weq3719));
    equaln #(12) e3720(.a(buffered_input), .b(12'b111010001000), .eq(weq3720));
    equaln #(12) e3721(.a(buffered_input), .b(12'b111010001001), .eq(weq3721));
    equaln #(12) e3722(.a(buffered_input), .b(12'b111010001010), .eq(weq3722));
    equaln #(12) e3723(.a(buffered_input), .b(12'b111010001011), .eq(weq3723));
    equaln #(12) e3724(.a(buffered_input), .b(12'b111010001100), .eq(weq3724));
    equaln #(12) e3725(.a(buffered_input), .b(12'b111010001101), .eq(weq3725));
    equaln #(12) e3726(.a(buffered_input), .b(12'b111010001110), .eq(weq3726));
    equaln #(12) e3727(.a(buffered_input), .b(12'b111010001111), .eq(weq3727));
    equaln #(12) e3728(.a(buffered_input), .b(12'b111010010000), .eq(weq3728));
    equaln #(12) e3729(.a(buffered_input), .b(12'b111010010001), .eq(weq3729));
    equaln #(12) e3730(.a(buffered_input), .b(12'b111010010010), .eq(weq3730));
    equaln #(12) e3731(.a(buffered_input), .b(12'b111010010011), .eq(weq3731));
    equaln #(12) e3732(.a(buffered_input), .b(12'b111010010100), .eq(weq3732));
    equaln #(12) e3733(.a(buffered_input), .b(12'b111010010101), .eq(weq3733));
    equaln #(12) e3734(.a(buffered_input), .b(12'b111010010110), .eq(weq3734));
    equaln #(12) e3735(.a(buffered_input), .b(12'b111010010111), .eq(weq3735));
    equaln #(12) e3736(.a(buffered_input), .b(12'b111010011000), .eq(weq3736));
    equaln #(12) e3737(.a(buffered_input), .b(12'b111010011001), .eq(weq3737));
    equaln #(12) e3738(.a(buffered_input), .b(12'b111010011010), .eq(weq3738));
    equaln #(12) e3739(.a(buffered_input), .b(12'b111010011011), .eq(weq3739));
    equaln #(12) e3740(.a(buffered_input), .b(12'b111010011100), .eq(weq3740));
    equaln #(12) e3741(.a(buffered_input), .b(12'b111010011101), .eq(weq3741));
    equaln #(12) e3742(.a(buffered_input), .b(12'b111010011110), .eq(weq3742));
    equaln #(12) e3743(.a(buffered_input), .b(12'b111010011111), .eq(weq3743));
    equaln #(12) e3744(.a(buffered_input), .b(12'b111010100000), .eq(weq3744));
    equaln #(12) e3745(.a(buffered_input), .b(12'b111010100001), .eq(weq3745));
    equaln #(12) e3746(.a(buffered_input), .b(12'b111010100010), .eq(weq3746));
    equaln #(12) e3747(.a(buffered_input), .b(12'b111010100011), .eq(weq3747));
    equaln #(12) e3748(.a(buffered_input), .b(12'b111010100100), .eq(weq3748));
    equaln #(12) e3749(.a(buffered_input), .b(12'b111010100101), .eq(weq3749));
    equaln #(12) e3750(.a(buffered_input), .b(12'b111010100110), .eq(weq3750));
    equaln #(12) e3751(.a(buffered_input), .b(12'b111010100111), .eq(weq3751));
    equaln #(12) e3752(.a(buffered_input), .b(12'b111010101000), .eq(weq3752));
    equaln #(12) e3753(.a(buffered_input), .b(12'b111010101001), .eq(weq3753));
    equaln #(12) e3754(.a(buffered_input), .b(12'b111010101010), .eq(weq3754));
    equaln #(12) e3755(.a(buffered_input), .b(12'b111010101011), .eq(weq3755));
    equaln #(12) e3756(.a(buffered_input), .b(12'b111010101100), .eq(weq3756));
    equaln #(12) e3757(.a(buffered_input), .b(12'b111010101101), .eq(weq3757));
    equaln #(12) e3758(.a(buffered_input), .b(12'b111010101110), .eq(weq3758));
    equaln #(12) e3759(.a(buffered_input), .b(12'b111010101111), .eq(weq3759));
    equaln #(12) e3760(.a(buffered_input), .b(12'b111010110000), .eq(weq3760));
    equaln #(12) e3761(.a(buffered_input), .b(12'b111010110001), .eq(weq3761));
    equaln #(12) e3762(.a(buffered_input), .b(12'b111010110010), .eq(weq3762));
    equaln #(12) e3763(.a(buffered_input), .b(12'b111010110011), .eq(weq3763));
    equaln #(12) e3764(.a(buffered_input), .b(12'b111010110100), .eq(weq3764));
    equaln #(12) e3765(.a(buffered_input), .b(12'b111010110101), .eq(weq3765));
    equaln #(12) e3766(.a(buffered_input), .b(12'b111010110110), .eq(weq3766));
    equaln #(12) e3767(.a(buffered_input), .b(12'b111010110111), .eq(weq3767));
    equaln #(12) e3768(.a(buffered_input), .b(12'b111010111000), .eq(weq3768));
    equaln #(12) e3769(.a(buffered_input), .b(12'b111010111001), .eq(weq3769));
    equaln #(12) e3770(.a(buffered_input), .b(12'b111010111010), .eq(weq3770));
    equaln #(12) e3771(.a(buffered_input), .b(12'b111010111011), .eq(weq3771));
    equaln #(12) e3772(.a(buffered_input), .b(12'b111010111100), .eq(weq3772));
    equaln #(12) e3773(.a(buffered_input), .b(12'b111010111101), .eq(weq3773));
    equaln #(12) e3774(.a(buffered_input), .b(12'b111010111110), .eq(weq3774));
    equaln #(12) e3775(.a(buffered_input), .b(12'b111010111111), .eq(weq3775));
    equaln #(12) e3776(.a(buffered_input), .b(12'b111011000000), .eq(weq3776));
    equaln #(12) e3777(.a(buffered_input), .b(12'b111011000001), .eq(weq3777));
    equaln #(12) e3778(.a(buffered_input), .b(12'b111011000010), .eq(weq3778));
    equaln #(12) e3779(.a(buffered_input), .b(12'b111011000011), .eq(weq3779));
    equaln #(12) e3780(.a(buffered_input), .b(12'b111011000100), .eq(weq3780));
    equaln #(12) e3781(.a(buffered_input), .b(12'b111011000101), .eq(weq3781));
    equaln #(12) e3782(.a(buffered_input), .b(12'b111011000110), .eq(weq3782));
    equaln #(12) e3783(.a(buffered_input), .b(12'b111011000111), .eq(weq3783));
    equaln #(12) e3784(.a(buffered_input), .b(12'b111011001000), .eq(weq3784));
    equaln #(12) e3785(.a(buffered_input), .b(12'b111011001001), .eq(weq3785));
    equaln #(12) e3786(.a(buffered_input), .b(12'b111011001010), .eq(weq3786));
    equaln #(12) e3787(.a(buffered_input), .b(12'b111011001011), .eq(weq3787));
    equaln #(12) e3788(.a(buffered_input), .b(12'b111011001100), .eq(weq3788));
    equaln #(12) e3789(.a(buffered_input), .b(12'b111011001101), .eq(weq3789));
    equaln #(12) e3790(.a(buffered_input), .b(12'b111011001110), .eq(weq3790));
    equaln #(12) e3791(.a(buffered_input), .b(12'b111011001111), .eq(weq3791));
    equaln #(12) e3792(.a(buffered_input), .b(12'b111011010000), .eq(weq3792));
    equaln #(12) e3793(.a(buffered_input), .b(12'b111011010001), .eq(weq3793));
    equaln #(12) e3794(.a(buffered_input), .b(12'b111011010010), .eq(weq3794));
    equaln #(12) e3795(.a(buffered_input), .b(12'b111011010011), .eq(weq3795));
    equaln #(12) e3796(.a(buffered_input), .b(12'b111011010100), .eq(weq3796));
    equaln #(12) e3797(.a(buffered_input), .b(12'b111011010101), .eq(weq3797));
    equaln #(12) e3798(.a(buffered_input), .b(12'b111011010110), .eq(weq3798));
    equaln #(12) e3799(.a(buffered_input), .b(12'b111011010111), .eq(weq3799));
    equaln #(12) e3800(.a(buffered_input), .b(12'b111011011000), .eq(weq3800));
    equaln #(12) e3801(.a(buffered_input), .b(12'b111011011001), .eq(weq3801));
    equaln #(12) e3802(.a(buffered_input), .b(12'b111011011010), .eq(weq3802));
    equaln #(12) e3803(.a(buffered_input), .b(12'b111011011011), .eq(weq3803));
    equaln #(12) e3804(.a(buffered_input), .b(12'b111011011100), .eq(weq3804));
    equaln #(12) e3805(.a(buffered_input), .b(12'b111011011101), .eq(weq3805));
    equaln #(12) e3806(.a(buffered_input), .b(12'b111011011110), .eq(weq3806));
    equaln #(12) e3807(.a(buffered_input), .b(12'b111011011111), .eq(weq3807));
    equaln #(12) e3808(.a(buffered_input), .b(12'b111011100000), .eq(weq3808));
    equaln #(12) e3809(.a(buffered_input), .b(12'b111011100001), .eq(weq3809));
    equaln #(12) e3810(.a(buffered_input), .b(12'b111011100010), .eq(weq3810));
    equaln #(12) e3811(.a(buffered_input), .b(12'b111011100011), .eq(weq3811));
    equaln #(12) e3812(.a(buffered_input), .b(12'b111011100100), .eq(weq3812));
    equaln #(12) e3813(.a(buffered_input), .b(12'b111011100101), .eq(weq3813));
    equaln #(12) e3814(.a(buffered_input), .b(12'b111011100110), .eq(weq3814));
    equaln #(12) e3815(.a(buffered_input), .b(12'b111011100111), .eq(weq3815));
    equaln #(12) e3816(.a(buffered_input), .b(12'b111011101000), .eq(weq3816));
    equaln #(12) e3817(.a(buffered_input), .b(12'b111011101001), .eq(weq3817));
    equaln #(12) e3818(.a(buffered_input), .b(12'b111011101010), .eq(weq3818));
    equaln #(12) e3819(.a(buffered_input), .b(12'b111011101011), .eq(weq3819));
    equaln #(12) e3820(.a(buffered_input), .b(12'b111011101100), .eq(weq3820));
    equaln #(12) e3821(.a(buffered_input), .b(12'b111011101101), .eq(weq3821));
    equaln #(12) e3822(.a(buffered_input), .b(12'b111011101110), .eq(weq3822));
    equaln #(12) e3823(.a(buffered_input), .b(12'b111011101111), .eq(weq3823));
    equaln #(12) e3824(.a(buffered_input), .b(12'b111011110000), .eq(weq3824));
    equaln #(12) e3825(.a(buffered_input), .b(12'b111011110001), .eq(weq3825));
    equaln #(12) e3826(.a(buffered_input), .b(12'b111011110010), .eq(weq3826));
    equaln #(12) e3827(.a(buffered_input), .b(12'b111011110011), .eq(weq3827));
    equaln #(12) e3828(.a(buffered_input), .b(12'b111011110100), .eq(weq3828));
    equaln #(12) e3829(.a(buffered_input), .b(12'b111011110101), .eq(weq3829));
    equaln #(12) e3830(.a(buffered_input), .b(12'b111011110110), .eq(weq3830));
    equaln #(12) e3831(.a(buffered_input), .b(12'b111011110111), .eq(weq3831));
    equaln #(12) e3832(.a(buffered_input), .b(12'b111011111000), .eq(weq3832));
    equaln #(12) e3833(.a(buffered_input), .b(12'b111011111001), .eq(weq3833));
    equaln #(12) e3834(.a(buffered_input), .b(12'b111011111010), .eq(weq3834));
    equaln #(12) e3835(.a(buffered_input), .b(12'b111011111011), .eq(weq3835));
    equaln #(12) e3836(.a(buffered_input), .b(12'b111011111100), .eq(weq3836));
    equaln #(12) e3837(.a(buffered_input), .b(12'b111011111101), .eq(weq3837));
    equaln #(12) e3838(.a(buffered_input), .b(12'b111011111110), .eq(weq3838));
    equaln #(12) e3839(.a(buffered_input), .b(12'b111011111111), .eq(weq3839));
    equaln #(12) e3840(.a(buffered_input), .b(12'b111100000000), .eq(weq3840));
    equaln #(12) e3841(.a(buffered_input), .b(12'b111100000001), .eq(weq3841));
    equaln #(12) e3842(.a(buffered_input), .b(12'b111100000010), .eq(weq3842));
    equaln #(12) e3843(.a(buffered_input), .b(12'b111100000011), .eq(weq3843));
    equaln #(12) e3844(.a(buffered_input), .b(12'b111100000100), .eq(weq3844));
    equaln #(12) e3845(.a(buffered_input), .b(12'b111100000101), .eq(weq3845));
    equaln #(12) e3846(.a(buffered_input), .b(12'b111100000110), .eq(weq3846));
    equaln #(12) e3847(.a(buffered_input), .b(12'b111100000111), .eq(weq3847));
    equaln #(12) e3848(.a(buffered_input), .b(12'b111100001000), .eq(weq3848));
    equaln #(12) e3849(.a(buffered_input), .b(12'b111100001001), .eq(weq3849));
    equaln #(12) e3850(.a(buffered_input), .b(12'b111100001010), .eq(weq3850));
    equaln #(12) e3851(.a(buffered_input), .b(12'b111100001011), .eq(weq3851));
    equaln #(12) e3852(.a(buffered_input), .b(12'b111100001100), .eq(weq3852));
    equaln #(12) e3853(.a(buffered_input), .b(12'b111100001101), .eq(weq3853));
    equaln #(12) e3854(.a(buffered_input), .b(12'b111100001110), .eq(weq3854));
    equaln #(12) e3855(.a(buffered_input), .b(12'b111100001111), .eq(weq3855));
    equaln #(12) e3856(.a(buffered_input), .b(12'b111100010000), .eq(weq3856));
    equaln #(12) e3857(.a(buffered_input), .b(12'b111100010001), .eq(weq3857));
    equaln #(12) e3858(.a(buffered_input), .b(12'b111100010010), .eq(weq3858));
    equaln #(12) e3859(.a(buffered_input), .b(12'b111100010011), .eq(weq3859));
    equaln #(12) e3860(.a(buffered_input), .b(12'b111100010100), .eq(weq3860));
    equaln #(12) e3861(.a(buffered_input), .b(12'b111100010101), .eq(weq3861));
    equaln #(12) e3862(.a(buffered_input), .b(12'b111100010110), .eq(weq3862));
    equaln #(12) e3863(.a(buffered_input), .b(12'b111100010111), .eq(weq3863));
    equaln #(12) e3864(.a(buffered_input), .b(12'b111100011000), .eq(weq3864));
    equaln #(12) e3865(.a(buffered_input), .b(12'b111100011001), .eq(weq3865));
    equaln #(12) e3866(.a(buffered_input), .b(12'b111100011010), .eq(weq3866));
    equaln #(12) e3867(.a(buffered_input), .b(12'b111100011011), .eq(weq3867));
    equaln #(12) e3868(.a(buffered_input), .b(12'b111100011100), .eq(weq3868));
    equaln #(12) e3869(.a(buffered_input), .b(12'b111100011101), .eq(weq3869));
    equaln #(12) e3870(.a(buffered_input), .b(12'b111100011110), .eq(weq3870));
    equaln #(12) e3871(.a(buffered_input), .b(12'b111100011111), .eq(weq3871));
    equaln #(12) e3872(.a(buffered_input), .b(12'b111100100000), .eq(weq3872));
    equaln #(12) e3873(.a(buffered_input), .b(12'b111100100001), .eq(weq3873));
    equaln #(12) e3874(.a(buffered_input), .b(12'b111100100010), .eq(weq3874));
    equaln #(12) e3875(.a(buffered_input), .b(12'b111100100011), .eq(weq3875));
    equaln #(12) e3876(.a(buffered_input), .b(12'b111100100100), .eq(weq3876));
    equaln #(12) e3877(.a(buffered_input), .b(12'b111100100101), .eq(weq3877));
    equaln #(12) e3878(.a(buffered_input), .b(12'b111100100110), .eq(weq3878));
    equaln #(12) e3879(.a(buffered_input), .b(12'b111100100111), .eq(weq3879));
    equaln #(12) e3880(.a(buffered_input), .b(12'b111100101000), .eq(weq3880));
    equaln #(12) e3881(.a(buffered_input), .b(12'b111100101001), .eq(weq3881));
    equaln #(12) e3882(.a(buffered_input), .b(12'b111100101010), .eq(weq3882));
    equaln #(12) e3883(.a(buffered_input), .b(12'b111100101011), .eq(weq3883));
    equaln #(12) e3884(.a(buffered_input), .b(12'b111100101100), .eq(weq3884));
    equaln #(12) e3885(.a(buffered_input), .b(12'b111100101101), .eq(weq3885));
    equaln #(12) e3886(.a(buffered_input), .b(12'b111100101110), .eq(weq3886));
    equaln #(12) e3887(.a(buffered_input), .b(12'b111100101111), .eq(weq3887));
    equaln #(12) e3888(.a(buffered_input), .b(12'b111100110000), .eq(weq3888));
    equaln #(12) e3889(.a(buffered_input), .b(12'b111100110001), .eq(weq3889));
    equaln #(12) e3890(.a(buffered_input), .b(12'b111100110010), .eq(weq3890));
    equaln #(12) e3891(.a(buffered_input), .b(12'b111100110011), .eq(weq3891));
    equaln #(12) e3892(.a(buffered_input), .b(12'b111100110100), .eq(weq3892));
    equaln #(12) e3893(.a(buffered_input), .b(12'b111100110101), .eq(weq3893));
    equaln #(12) e3894(.a(buffered_input), .b(12'b111100110110), .eq(weq3894));
    equaln #(12) e3895(.a(buffered_input), .b(12'b111100110111), .eq(weq3895));
    equaln #(12) e3896(.a(buffered_input), .b(12'b111100111000), .eq(weq3896));
    equaln #(12) e3897(.a(buffered_input), .b(12'b111100111001), .eq(weq3897));
    equaln #(12) e3898(.a(buffered_input), .b(12'b111100111010), .eq(weq3898));
    equaln #(12) e3899(.a(buffered_input), .b(12'b111100111011), .eq(weq3899));
    equaln #(12) e3900(.a(buffered_input), .b(12'b111100111100), .eq(weq3900));
    equaln #(12) e3901(.a(buffered_input), .b(12'b111100111101), .eq(weq3901));
    equaln #(12) e3902(.a(buffered_input), .b(12'b111100111110), .eq(weq3902));
    equaln #(12) e3903(.a(buffered_input), .b(12'b111100111111), .eq(weq3903));
    equaln #(12) e3904(.a(buffered_input), .b(12'b111101000000), .eq(weq3904));
    equaln #(12) e3905(.a(buffered_input), .b(12'b111101000001), .eq(weq3905));
    equaln #(12) e3906(.a(buffered_input), .b(12'b111101000010), .eq(weq3906));
    equaln #(12) e3907(.a(buffered_input), .b(12'b111101000011), .eq(weq3907));
    equaln #(12) e3908(.a(buffered_input), .b(12'b111101000100), .eq(weq3908));
    equaln #(12) e3909(.a(buffered_input), .b(12'b111101000101), .eq(weq3909));
    equaln #(12) e3910(.a(buffered_input), .b(12'b111101000110), .eq(weq3910));
    equaln #(12) e3911(.a(buffered_input), .b(12'b111101000111), .eq(weq3911));
    equaln #(12) e3912(.a(buffered_input), .b(12'b111101001000), .eq(weq3912));
    equaln #(12) e3913(.a(buffered_input), .b(12'b111101001001), .eq(weq3913));
    equaln #(12) e3914(.a(buffered_input), .b(12'b111101001010), .eq(weq3914));
    equaln #(12) e3915(.a(buffered_input), .b(12'b111101001011), .eq(weq3915));
    equaln #(12) e3916(.a(buffered_input), .b(12'b111101001100), .eq(weq3916));
    equaln #(12) e3917(.a(buffered_input), .b(12'b111101001101), .eq(weq3917));
    equaln #(12) e3918(.a(buffered_input), .b(12'b111101001110), .eq(weq3918));
    equaln #(12) e3919(.a(buffered_input), .b(12'b111101001111), .eq(weq3919));
    equaln #(12) e3920(.a(buffered_input), .b(12'b111101010000), .eq(weq3920));
    equaln #(12) e3921(.a(buffered_input), .b(12'b111101010001), .eq(weq3921));
    equaln #(12) e3922(.a(buffered_input), .b(12'b111101010010), .eq(weq3922));
    equaln #(12) e3923(.a(buffered_input), .b(12'b111101010011), .eq(weq3923));
    equaln #(12) e3924(.a(buffered_input), .b(12'b111101010100), .eq(weq3924));
    equaln #(12) e3925(.a(buffered_input), .b(12'b111101010101), .eq(weq3925));
    equaln #(12) e3926(.a(buffered_input), .b(12'b111101010110), .eq(weq3926));
    equaln #(12) e3927(.a(buffered_input), .b(12'b111101010111), .eq(weq3927));
    equaln #(12) e3928(.a(buffered_input), .b(12'b111101011000), .eq(weq3928));
    equaln #(12) e3929(.a(buffered_input), .b(12'b111101011001), .eq(weq3929));
    equaln #(12) e3930(.a(buffered_input), .b(12'b111101011010), .eq(weq3930));
    equaln #(12) e3931(.a(buffered_input), .b(12'b111101011011), .eq(weq3931));
    equaln #(12) e3932(.a(buffered_input), .b(12'b111101011100), .eq(weq3932));
    equaln #(12) e3933(.a(buffered_input), .b(12'b111101011101), .eq(weq3933));
    equaln #(12) e3934(.a(buffered_input), .b(12'b111101011110), .eq(weq3934));
    equaln #(12) e3935(.a(buffered_input), .b(12'b111101011111), .eq(weq3935));
    equaln #(12) e3936(.a(buffered_input), .b(12'b111101100000), .eq(weq3936));
    equaln #(12) e3937(.a(buffered_input), .b(12'b111101100001), .eq(weq3937));
    equaln #(12) e3938(.a(buffered_input), .b(12'b111101100010), .eq(weq3938));
    equaln #(12) e3939(.a(buffered_input), .b(12'b111101100011), .eq(weq3939));
    equaln #(12) e3940(.a(buffered_input), .b(12'b111101100100), .eq(weq3940));
    equaln #(12) e3941(.a(buffered_input), .b(12'b111101100101), .eq(weq3941));
    equaln #(12) e3942(.a(buffered_input), .b(12'b111101100110), .eq(weq3942));
    equaln #(12) e3943(.a(buffered_input), .b(12'b111101100111), .eq(weq3943));
    equaln #(12) e3944(.a(buffered_input), .b(12'b111101101000), .eq(weq3944));
    equaln #(12) e3945(.a(buffered_input), .b(12'b111101101001), .eq(weq3945));
    equaln #(12) e3946(.a(buffered_input), .b(12'b111101101010), .eq(weq3946));
    equaln #(12) e3947(.a(buffered_input), .b(12'b111101101011), .eq(weq3947));
    equaln #(12) e3948(.a(buffered_input), .b(12'b111101101100), .eq(weq3948));
    equaln #(12) e3949(.a(buffered_input), .b(12'b111101101101), .eq(weq3949));
    equaln #(12) e3950(.a(buffered_input), .b(12'b111101101110), .eq(weq3950));
    equaln #(12) e3951(.a(buffered_input), .b(12'b111101101111), .eq(weq3951));
    equaln #(12) e3952(.a(buffered_input), .b(12'b111101110000), .eq(weq3952));
    equaln #(12) e3953(.a(buffered_input), .b(12'b111101110001), .eq(weq3953));
    equaln #(12) e3954(.a(buffered_input), .b(12'b111101110010), .eq(weq3954));
    equaln #(12) e3955(.a(buffered_input), .b(12'b111101110011), .eq(weq3955));
    equaln #(12) e3956(.a(buffered_input), .b(12'b111101110100), .eq(weq3956));
    equaln #(12) e3957(.a(buffered_input), .b(12'b111101110101), .eq(weq3957));
    equaln #(12) e3958(.a(buffered_input), .b(12'b111101110110), .eq(weq3958));
    equaln #(12) e3959(.a(buffered_input), .b(12'b111101110111), .eq(weq3959));
    equaln #(12) e3960(.a(buffered_input), .b(12'b111101111000), .eq(weq3960));
    equaln #(12) e3961(.a(buffered_input), .b(12'b111101111001), .eq(weq3961));
    equaln #(12) e3962(.a(buffered_input), .b(12'b111101111010), .eq(weq3962));
    equaln #(12) e3963(.a(buffered_input), .b(12'b111101111011), .eq(weq3963));
    equaln #(12) e3964(.a(buffered_input), .b(12'b111101111100), .eq(weq3964));
    equaln #(12) e3965(.a(buffered_input), .b(12'b111101111101), .eq(weq3965));
    equaln #(12) e3966(.a(buffered_input), .b(12'b111101111110), .eq(weq3966));
    equaln #(12) e3967(.a(buffered_input), .b(12'b111101111111), .eq(weq3967));
    equaln #(12) e3968(.a(buffered_input), .b(12'b111110000000), .eq(weq3968));
    equaln #(12) e3969(.a(buffered_input), .b(12'b111110000001), .eq(weq3969));
    equaln #(12) e3970(.a(buffered_input), .b(12'b111110000010), .eq(weq3970));
    equaln #(12) e3971(.a(buffered_input), .b(12'b111110000011), .eq(weq3971));
    equaln #(12) e3972(.a(buffered_input), .b(12'b111110000100), .eq(weq3972));
    equaln #(12) e3973(.a(buffered_input), .b(12'b111110000101), .eq(weq3973));
    equaln #(12) e3974(.a(buffered_input), .b(12'b111110000110), .eq(weq3974));
    equaln #(12) e3975(.a(buffered_input), .b(12'b111110000111), .eq(weq3975));
    equaln #(12) e3976(.a(buffered_input), .b(12'b111110001000), .eq(weq3976));
    equaln #(12) e3977(.a(buffered_input), .b(12'b111110001001), .eq(weq3977));
    equaln #(12) e3978(.a(buffered_input), .b(12'b111110001010), .eq(weq3978));
    equaln #(12) e3979(.a(buffered_input), .b(12'b111110001011), .eq(weq3979));
    equaln #(12) e3980(.a(buffered_input), .b(12'b111110001100), .eq(weq3980));
    equaln #(12) e3981(.a(buffered_input), .b(12'b111110001101), .eq(weq3981));
    equaln #(12) e3982(.a(buffered_input), .b(12'b111110001110), .eq(weq3982));
    equaln #(12) e3983(.a(buffered_input), .b(12'b111110001111), .eq(weq3983));
    equaln #(12) e3984(.a(buffered_input), .b(12'b111110010000), .eq(weq3984));
    equaln #(12) e3985(.a(buffered_input), .b(12'b111110010001), .eq(weq3985));
    equaln #(12) e3986(.a(buffered_input), .b(12'b111110010010), .eq(weq3986));
    equaln #(12) e3987(.a(buffered_input), .b(12'b111110010011), .eq(weq3987));
    equaln #(12) e3988(.a(buffered_input), .b(12'b111110010100), .eq(weq3988));
    equaln #(12) e3989(.a(buffered_input), .b(12'b111110010101), .eq(weq3989));
    equaln #(12) e3990(.a(buffered_input), .b(12'b111110010110), .eq(weq3990));
    equaln #(12) e3991(.a(buffered_input), .b(12'b111110010111), .eq(weq3991));
    equaln #(12) e3992(.a(buffered_input), .b(12'b111110011000), .eq(weq3992));
    equaln #(12) e3993(.a(buffered_input), .b(12'b111110011001), .eq(weq3993));
    equaln #(12) e3994(.a(buffered_input), .b(12'b111110011010), .eq(weq3994));
    equaln #(12) e3995(.a(buffered_input), .b(12'b111110011011), .eq(weq3995));
    equaln #(12) e3996(.a(buffered_input), .b(12'b111110011100), .eq(weq3996));
    equaln #(12) e3997(.a(buffered_input), .b(12'b111110011101), .eq(weq3997));
    equaln #(12) e3998(.a(buffered_input), .b(12'b111110011110), .eq(weq3998));
    equaln #(12) e3999(.a(buffered_input), .b(12'b111110011111), .eq(weq3999));
    equaln #(12) e4000(.a(buffered_input), .b(12'b111110100000), .eq(weq4000));
    equaln #(12) e4001(.a(buffered_input), .b(12'b111110100001), .eq(weq4001));
    equaln #(12) e4002(.a(buffered_input), .b(12'b111110100010), .eq(weq4002));
    equaln #(12) e4003(.a(buffered_input), .b(12'b111110100011), .eq(weq4003));
    equaln #(12) e4004(.a(buffered_input), .b(12'b111110100100), .eq(weq4004));
    equaln #(12) e4005(.a(buffered_input), .b(12'b111110100101), .eq(weq4005));
    equaln #(12) e4006(.a(buffered_input), .b(12'b111110100110), .eq(weq4006));
    equaln #(12) e4007(.a(buffered_input), .b(12'b111110100111), .eq(weq4007));
    equaln #(12) e4008(.a(buffered_input), .b(12'b111110101000), .eq(weq4008));
    equaln #(12) e4009(.a(buffered_input), .b(12'b111110101001), .eq(weq4009));
    equaln #(12) e4010(.a(buffered_input), .b(12'b111110101010), .eq(weq4010));
    equaln #(12) e4011(.a(buffered_input), .b(12'b111110101011), .eq(weq4011));
    equaln #(12) e4012(.a(buffered_input), .b(12'b111110101100), .eq(weq4012));
    equaln #(12) e4013(.a(buffered_input), .b(12'b111110101101), .eq(weq4013));
    equaln #(12) e4014(.a(buffered_input), .b(12'b111110101110), .eq(weq4014));
    equaln #(12) e4015(.a(buffered_input), .b(12'b111110101111), .eq(weq4015));
    equaln #(12) e4016(.a(buffered_input), .b(12'b111110110000), .eq(weq4016));
    equaln #(12) e4017(.a(buffered_input), .b(12'b111110110001), .eq(weq4017));
    equaln #(12) e4018(.a(buffered_input), .b(12'b111110110010), .eq(weq4018));
    equaln #(12) e4019(.a(buffered_input), .b(12'b111110110011), .eq(weq4019));
    equaln #(12) e4020(.a(buffered_input), .b(12'b111110110100), .eq(weq4020));
    equaln #(12) e4021(.a(buffered_input), .b(12'b111110110101), .eq(weq4021));
    equaln #(12) e4022(.a(buffered_input), .b(12'b111110110110), .eq(weq4022));
    equaln #(12) e4023(.a(buffered_input), .b(12'b111110110111), .eq(weq4023));
    equaln #(12) e4024(.a(buffered_input), .b(12'b111110111000), .eq(weq4024));
    equaln #(12) e4025(.a(buffered_input), .b(12'b111110111001), .eq(weq4025));
    equaln #(12) e4026(.a(buffered_input), .b(12'b111110111010), .eq(weq4026));
    equaln #(12) e4027(.a(buffered_input), .b(12'b111110111011), .eq(weq4027));
    equaln #(12) e4028(.a(buffered_input), .b(12'b111110111100), .eq(weq4028));
    equaln #(12) e4029(.a(buffered_input), .b(12'b111110111101), .eq(weq4029));
    equaln #(12) e4030(.a(buffered_input), .b(12'b111110111110), .eq(weq4030));
    equaln #(12) e4031(.a(buffered_input), .b(12'b111110111111), .eq(weq4031));
    equaln #(12) e4032(.a(buffered_input), .b(12'b111111000000), .eq(weq4032));
    equaln #(12) e4033(.a(buffered_input), .b(12'b111111000001), .eq(weq4033));
    equaln #(12) e4034(.a(buffered_input), .b(12'b111111000010), .eq(weq4034));
    equaln #(12) e4035(.a(buffered_input), .b(12'b111111000011), .eq(weq4035));
    equaln #(12) e4036(.a(buffered_input), .b(12'b111111000100), .eq(weq4036));
    equaln #(12) e4037(.a(buffered_input), .b(12'b111111000101), .eq(weq4037));
    equaln #(12) e4038(.a(buffered_input), .b(12'b111111000110), .eq(weq4038));
    equaln #(12) e4039(.a(buffered_input), .b(12'b111111000111), .eq(weq4039));
    equaln #(12) e4040(.a(buffered_input), .b(12'b111111001000), .eq(weq4040));
    equaln #(12) e4041(.a(buffered_input), .b(12'b111111001001), .eq(weq4041));
    equaln #(12) e4042(.a(buffered_input), .b(12'b111111001010), .eq(weq4042));
    equaln #(12) e4043(.a(buffered_input), .b(12'b111111001011), .eq(weq4043));
    equaln #(12) e4044(.a(buffered_input), .b(12'b111111001100), .eq(weq4044));
    equaln #(12) e4045(.a(buffered_input), .b(12'b111111001101), .eq(weq4045));
    equaln #(12) e4046(.a(buffered_input), .b(12'b111111001110), .eq(weq4046));
    equaln #(12) e4047(.a(buffered_input), .b(12'b111111001111), .eq(weq4047));
    equaln #(12) e4048(.a(buffered_input), .b(12'b111111010000), .eq(weq4048));
    equaln #(12) e4049(.a(buffered_input), .b(12'b111111010001), .eq(weq4049));
    equaln #(12) e4050(.a(buffered_input), .b(12'b111111010010), .eq(weq4050));
    equaln #(12) e4051(.a(buffered_input), .b(12'b111111010011), .eq(weq4051));
    equaln #(12) e4052(.a(buffered_input), .b(12'b111111010100), .eq(weq4052));
    equaln #(12) e4053(.a(buffered_input), .b(12'b111111010101), .eq(weq4053));
    equaln #(12) e4054(.a(buffered_input), .b(12'b111111010110), .eq(weq4054));
    equaln #(12) e4055(.a(buffered_input), .b(12'b111111010111), .eq(weq4055));
    equaln #(12) e4056(.a(buffered_input), .b(12'b111111011000), .eq(weq4056));
    equaln #(12) e4057(.a(buffered_input), .b(12'b111111011001), .eq(weq4057));
    equaln #(12) e4058(.a(buffered_input), .b(12'b111111011010), .eq(weq4058));
    equaln #(12) e4059(.a(buffered_input), .b(12'b111111011011), .eq(weq4059));
    equaln #(12) e4060(.a(buffered_input), .b(12'b111111011100), .eq(weq4060));
    equaln #(12) e4061(.a(buffered_input), .b(12'b111111011101), .eq(weq4061));
    equaln #(12) e4062(.a(buffered_input), .b(12'b111111011110), .eq(weq4062));
    equaln #(12) e4063(.a(buffered_input), .b(12'b111111011111), .eq(weq4063));
    equaln #(12) e4064(.a(buffered_input), .b(12'b111111100000), .eq(weq4064));
    equaln #(12) e4065(.a(buffered_input), .b(12'b111111100001), .eq(weq4065));
    equaln #(12) e4066(.a(buffered_input), .b(12'b111111100010), .eq(weq4066));
    equaln #(12) e4067(.a(buffered_input), .b(12'b111111100011), .eq(weq4067));
    equaln #(12) e4068(.a(buffered_input), .b(12'b111111100100), .eq(weq4068));
    equaln #(12) e4069(.a(buffered_input), .b(12'b111111100101), .eq(weq4069));
    equaln #(12) e4070(.a(buffered_input), .b(12'b111111100110), .eq(weq4070));
    equaln #(12) e4071(.a(buffered_input), .b(12'b111111100111), .eq(weq4071));
    equaln #(12) e4072(.a(buffered_input), .b(12'b111111101000), .eq(weq4072));
    equaln #(12) e4073(.a(buffered_input), .b(12'b111111101001), .eq(weq4073));
    equaln #(12) e4074(.a(buffered_input), .b(12'b111111101010), .eq(weq4074));
    equaln #(12) e4075(.a(buffered_input), .b(12'b111111101011), .eq(weq4075));
    equaln #(12) e4076(.a(buffered_input), .b(12'b111111101100), .eq(weq4076));
    equaln #(12) e4077(.a(buffered_input), .b(12'b111111101101), .eq(weq4077));
    equaln #(12) e4078(.a(buffered_input), .b(12'b111111101110), .eq(weq4078));
    equaln #(12) e4079(.a(buffered_input), .b(12'b111111101111), .eq(weq4079));
    equaln #(12) e4080(.a(buffered_input), .b(12'b111111110000), .eq(weq4080));
    equaln #(12) e4081(.a(buffered_input), .b(12'b111111110001), .eq(weq4081));
    equaln #(12) e4082(.a(buffered_input), .b(12'b111111110010), .eq(weq4082));
    equaln #(12) e4083(.a(buffered_input), .b(12'b111111110011), .eq(weq4083));
    equaln #(12) e4084(.a(buffered_input), .b(12'b111111110100), .eq(weq4084));
    equaln #(12) e4085(.a(buffered_input), .b(12'b111111110101), .eq(weq4085));
    equaln #(12) e4086(.a(buffered_input), .b(12'b111111110110), .eq(weq4086));
    equaln #(12) e4087(.a(buffered_input), .b(12'b111111110111), .eq(weq4087));
    equaln #(12) e4088(.a(buffered_input), .b(12'b111111111000), .eq(weq4088));
    equaln #(12) e4089(.a(buffered_input), .b(12'b111111111001), .eq(weq4089));
    equaln #(12) e4090(.a(buffered_input), .b(12'b111111111010), .eq(weq4090));
    equaln #(12) e4091(.a(buffered_input), .b(12'b111111111011), .eq(weq4091));
    equaln #(12) e4092(.a(buffered_input), .b(12'b111111111100), .eq(weq4092));
    equaln #(12) e4093(.a(buffered_input), .b(12'b111111111101), .eq(weq4093));
    equaln #(12) e4094(.a(buffered_input), .b(12'b111111111110), .eq(weq4094));
    equaln #(12) e4095(.a(buffered_input), .b(12'b111111111111), .eq(weq4095));


    wire [4095:0] weq_concat;
    assign weq_concat = {weq4095, weq4094, weq4093, weq4092, weq4091, weq4090, weq4089, weq4088, weq4087, weq4086, weq4085, weq4084, weq4083, weq4082, weq4081, weq4080, weq4079, weq4078, weq4077, weq4076, weq4075, weq4074, weq4073, weq4072, weq4071, weq4070, weq4069, weq4068, weq4067, weq4066, weq4065, weq4064, weq4063, weq4062, weq4061, weq4060, weq4059, weq4058, weq4057, weq4056, weq4055, weq4054, weq4053, weq4052, weq4051, weq4050, weq4049, weq4048, weq4047, weq4046, weq4045, weq4044, weq4043, weq4042, weq4041, weq4040, weq4039, weq4038, weq4037, weq4036, weq4035, weq4034, weq4033, weq4032, weq4031, weq4030, weq4029, weq4028, weq4027, weq4026, weq4025, weq4024, weq4023, weq4022, weq4021, weq4020, weq4019, weq4018, weq4017, weq4016, weq4015, weq4014, weq4013, weq4012, weq4011, weq4010, weq4009, weq4008, weq4007, weq4006, weq4005, weq4004, weq4003, weq4002, weq4001, weq4000, weq3999, weq3998, weq3997, weq3996, weq3995, weq3994, weq3993, weq3992, weq3991, weq3990, weq3989, weq3988, weq3987, weq3986, weq3985, weq3984, weq3983, weq3982, weq3981, weq3980, weq3979, weq3978, weq3977, weq3976, weq3975, weq3974, weq3973, weq3972, weq3971, weq3970, weq3969, weq3968, weq3967, weq3966, weq3965, weq3964, weq3963, weq3962, weq3961, weq3960, weq3959, weq3958, weq3957, weq3956, weq3955, weq3954, weq3953, weq3952, weq3951, weq3950, weq3949, weq3948, weq3947, weq3946, weq3945, weq3944, weq3943, weq3942, weq3941, weq3940, weq3939, weq3938, weq3937, weq3936, weq3935, weq3934, weq3933, weq3932, weq3931, weq3930, weq3929, weq3928, weq3927, weq3926, weq3925, weq3924, weq3923, weq3922, weq3921, weq3920, weq3919, weq3918, weq3917, weq3916, weq3915, weq3914, weq3913, weq3912, weq3911, weq3910, weq3909, weq3908, weq3907, weq3906, weq3905, weq3904, weq3903, weq3902, weq3901, weq3900, weq3899, weq3898, weq3897, weq3896, weq3895, weq3894, weq3893, weq3892, weq3891, weq3890, weq3889, weq3888, weq3887, weq3886, weq3885, weq3884, weq3883, weq3882, weq3881, weq3880, weq3879, weq3878, weq3877, weq3876, weq3875, weq3874, weq3873, weq3872, weq3871, weq3870, weq3869, weq3868, weq3867, weq3866, weq3865, weq3864, weq3863, weq3862, weq3861, weq3860, weq3859, weq3858, weq3857, weq3856, weq3855, weq3854, weq3853, weq3852, weq3851, weq3850, weq3849, weq3848, weq3847, weq3846, weq3845, weq3844, weq3843, weq3842, weq3841, weq3840, weq3839, weq3838, weq3837, weq3836, weq3835, weq3834, weq3833, weq3832, weq3831, weq3830, weq3829, weq3828, weq3827, weq3826, weq3825, weq3824, weq3823, weq3822, weq3821, weq3820, weq3819, weq3818, weq3817, weq3816, weq3815, weq3814, weq3813, weq3812, weq3811, weq3810, weq3809, weq3808, weq3807, weq3806, weq3805, weq3804, weq3803, weq3802, weq3801, weq3800, weq3799, weq3798, weq3797, weq3796, weq3795, weq3794, weq3793, weq3792, weq3791, weq3790, weq3789, weq3788, weq3787, weq3786, weq3785, weq3784, weq3783, weq3782, weq3781, weq3780, weq3779, weq3778, weq3777, weq3776, weq3775, weq3774, weq3773, weq3772, weq3771, weq3770, weq3769, weq3768, weq3767, weq3766, weq3765, weq3764, weq3763, weq3762, weq3761, weq3760, weq3759, weq3758, weq3757, weq3756, weq3755, weq3754, weq3753, weq3752, weq3751, weq3750, weq3749, weq3748, weq3747, weq3746, weq3745, weq3744, weq3743, weq3742, weq3741, weq3740, weq3739, weq3738, weq3737, weq3736, weq3735, weq3734, weq3733, weq3732, weq3731, weq3730, weq3729, weq3728, weq3727, weq3726, weq3725, weq3724, weq3723, weq3722, weq3721, weq3720, weq3719, weq3718, weq3717, weq3716, weq3715, weq3714, weq3713, weq3712, weq3711, weq3710, weq3709, weq3708, weq3707, weq3706, weq3705, weq3704, weq3703, weq3702, weq3701, weq3700, weq3699, weq3698, weq3697, weq3696, weq3695, weq3694, weq3693, weq3692, weq3691, weq3690, weq3689, weq3688, weq3687, weq3686, weq3685, weq3684, weq3683, weq3682, weq3681, weq3680, weq3679, weq3678, weq3677, weq3676, weq3675, weq3674, weq3673, weq3672, weq3671, weq3670, weq3669, weq3668, weq3667, weq3666, weq3665, weq3664, weq3663, weq3662, weq3661, weq3660, weq3659, weq3658, weq3657, weq3656, weq3655, weq3654, weq3653, weq3652, weq3651, weq3650, weq3649, weq3648, weq3647, weq3646, weq3645, weq3644, weq3643, weq3642, weq3641, weq3640, weq3639, weq3638, weq3637, weq3636, weq3635, weq3634, weq3633, weq3632, weq3631, weq3630, weq3629, weq3628, weq3627, weq3626, weq3625, weq3624, weq3623, weq3622, weq3621, weq3620, weq3619, weq3618, weq3617, weq3616, weq3615, weq3614, weq3613, weq3612, weq3611, weq3610, weq3609, weq3608, weq3607, weq3606, weq3605, weq3604, weq3603, weq3602, weq3601, weq3600, weq3599, weq3598, weq3597, weq3596, weq3595, weq3594, weq3593, weq3592, weq3591, weq3590, weq3589, weq3588, weq3587, weq3586, weq3585, weq3584, weq3583, weq3582, weq3581, weq3580, weq3579, weq3578, weq3577, weq3576, weq3575, weq3574, weq3573, weq3572, weq3571, weq3570, weq3569, weq3568, weq3567, weq3566, weq3565, weq3564, weq3563, weq3562, weq3561, weq3560, weq3559, weq3558, weq3557, weq3556, weq3555, weq3554, weq3553, weq3552, weq3551, weq3550, weq3549, weq3548, weq3547, weq3546, weq3545, weq3544, weq3543, weq3542, weq3541, weq3540, weq3539, weq3538, weq3537, weq3536, weq3535, weq3534, weq3533, weq3532, weq3531, weq3530, weq3529, weq3528, weq3527, weq3526, weq3525, weq3524, weq3523, weq3522, weq3521, weq3520, weq3519, weq3518, weq3517, weq3516, weq3515, weq3514, weq3513, weq3512, weq3511, weq3510, weq3509, weq3508, weq3507, weq3506, weq3505, weq3504, weq3503, weq3502, weq3501, weq3500, weq3499, weq3498, weq3497, weq3496, weq3495, weq3494, weq3493, weq3492, weq3491, weq3490, weq3489, weq3488, weq3487, weq3486, weq3485, weq3484, weq3483, weq3482, weq3481, weq3480, weq3479, weq3478, weq3477, weq3476, weq3475, weq3474, weq3473, weq3472, weq3471, weq3470, weq3469, weq3468, weq3467, weq3466, weq3465, weq3464, weq3463, weq3462, weq3461, weq3460, weq3459, weq3458, weq3457, weq3456, weq3455, weq3454, weq3453, weq3452, weq3451, weq3450, weq3449, weq3448, weq3447, weq3446, weq3445, weq3444, weq3443, weq3442, weq3441, weq3440, weq3439, weq3438, weq3437, weq3436, weq3435, weq3434, weq3433, weq3432, weq3431, weq3430, weq3429, weq3428, weq3427, weq3426, weq3425, weq3424, weq3423, weq3422, weq3421, weq3420, weq3419, weq3418, weq3417, weq3416, weq3415, weq3414, weq3413, weq3412, weq3411, weq3410, weq3409, weq3408, weq3407, weq3406, weq3405, weq3404, weq3403, weq3402, weq3401, weq3400, weq3399, weq3398, weq3397, weq3396, weq3395, weq3394, weq3393, weq3392, weq3391, weq3390, weq3389, weq3388, weq3387, weq3386, weq3385, weq3384, weq3383, weq3382, weq3381, weq3380, weq3379, weq3378, weq3377, weq3376, weq3375, weq3374, weq3373, weq3372, weq3371, weq3370, weq3369, weq3368, weq3367, weq3366, weq3365, weq3364, weq3363, weq3362, weq3361, weq3360, weq3359, weq3358, weq3357, weq3356, weq3355, weq3354, weq3353, weq3352, weq3351, weq3350, weq3349, weq3348, weq3347, weq3346, weq3345, weq3344, weq3343, weq3342, weq3341, weq3340, weq3339, weq3338, weq3337, weq3336, weq3335, weq3334, weq3333, weq3332, weq3331, weq3330, weq3329, weq3328, weq3327, weq3326, weq3325, weq3324, weq3323, weq3322, weq3321, weq3320, weq3319, weq3318, weq3317, weq3316, weq3315, weq3314, weq3313, weq3312, weq3311, weq3310, weq3309, weq3308, weq3307, weq3306, weq3305, weq3304, weq3303, weq3302, weq3301, weq3300, weq3299, weq3298, weq3297, weq3296, weq3295, weq3294, weq3293, weq3292, weq3291, weq3290, weq3289, weq3288, weq3287, weq3286, weq3285, weq3284, weq3283, weq3282, weq3281, weq3280, weq3279, weq3278, weq3277, weq3276, weq3275, weq3274, weq3273, weq3272, weq3271, weq3270, weq3269, weq3268, weq3267, weq3266, weq3265, weq3264, weq3263, weq3262, weq3261, weq3260, weq3259, weq3258, weq3257, weq3256, weq3255, weq3254, weq3253, weq3252, weq3251, weq3250, weq3249, weq3248, weq3247, weq3246, weq3245, weq3244, weq3243, weq3242, weq3241, weq3240, weq3239, weq3238, weq3237, weq3236, weq3235, weq3234, weq3233, weq3232, weq3231, weq3230, weq3229, weq3228, weq3227, weq3226, weq3225, weq3224, weq3223, weq3222, weq3221, weq3220, weq3219, weq3218, weq3217, weq3216, weq3215, weq3214, weq3213, weq3212, weq3211, weq3210, weq3209, weq3208, weq3207, weq3206, weq3205, weq3204, weq3203, weq3202, weq3201, weq3200, weq3199, weq3198, weq3197, weq3196, weq3195, weq3194, weq3193, weq3192, weq3191, weq3190, weq3189, weq3188, weq3187, weq3186, weq3185, weq3184, weq3183, weq3182, weq3181, weq3180, weq3179, weq3178, weq3177, weq3176, weq3175, weq3174, weq3173, weq3172, weq3171, weq3170, weq3169, weq3168, weq3167, weq3166, weq3165, weq3164, weq3163, weq3162, weq3161, weq3160, weq3159, weq3158, weq3157, weq3156, weq3155, weq3154, weq3153, weq3152, weq3151, weq3150, weq3149, weq3148, weq3147, weq3146, weq3145, weq3144, weq3143, weq3142, weq3141, weq3140, weq3139, weq3138, weq3137, weq3136, weq3135, weq3134, weq3133, weq3132, weq3131, weq3130, weq3129, weq3128, weq3127, weq3126, weq3125, weq3124, weq3123, weq3122, weq3121, weq3120, weq3119, weq3118, weq3117, weq3116, weq3115, weq3114, weq3113, weq3112, weq3111, weq3110, weq3109, weq3108, weq3107, weq3106, weq3105, weq3104, weq3103, weq3102, weq3101, weq3100, weq3099, weq3098, weq3097, weq3096, weq3095, weq3094, weq3093, weq3092, weq3091, weq3090, weq3089, weq3088, weq3087, weq3086, weq3085, weq3084, weq3083, weq3082, weq3081, weq3080, weq3079, weq3078, weq3077, weq3076, weq3075, weq3074, weq3073, weq3072, weq3071, weq3070, weq3069, weq3068, weq3067, weq3066, weq3065, weq3064, weq3063, weq3062, weq3061, weq3060, weq3059, weq3058, weq3057, weq3056, weq3055, weq3054, weq3053, weq3052, weq3051, weq3050, weq3049, weq3048, weq3047, weq3046, weq3045, weq3044, weq3043, weq3042, weq3041, weq3040, weq3039, weq3038, weq3037, weq3036, weq3035, weq3034, weq3033, weq3032, weq3031, weq3030, weq3029, weq3028, weq3027, weq3026, weq3025, weq3024, weq3023, weq3022, weq3021, weq3020, weq3019, weq3018, weq3017, weq3016, weq3015, weq3014, weq3013, weq3012, weq3011, weq3010, weq3009, weq3008, weq3007, weq3006, weq3005, weq3004, weq3003, weq3002, weq3001, weq3000, weq2999, weq2998, weq2997, weq2996, weq2995, weq2994, weq2993, weq2992, weq2991, weq2990, weq2989, weq2988, weq2987, weq2986, weq2985, weq2984, weq2983, weq2982, weq2981, weq2980, weq2979, weq2978, weq2977, weq2976, weq2975, weq2974, weq2973, weq2972, weq2971, weq2970, weq2969, weq2968, weq2967, weq2966, weq2965, weq2964, weq2963, weq2962, weq2961, weq2960, weq2959, weq2958, weq2957, weq2956, weq2955, weq2954, weq2953, weq2952, weq2951, weq2950, weq2949, weq2948, weq2947, weq2946, weq2945, weq2944, weq2943, weq2942, weq2941, weq2940, weq2939, weq2938, weq2937, weq2936, weq2935, weq2934, weq2933, weq2932, weq2931, weq2930, weq2929, weq2928, weq2927, weq2926, weq2925, weq2924, weq2923, weq2922, weq2921, weq2920, weq2919, weq2918, weq2917, weq2916, weq2915, weq2914, weq2913, weq2912, weq2911, weq2910, weq2909, weq2908, weq2907, weq2906, weq2905, weq2904, weq2903, weq2902, weq2901, weq2900, weq2899, weq2898, weq2897, weq2896, weq2895, weq2894, weq2893, weq2892, weq2891, weq2890, weq2889, weq2888, weq2887, weq2886, weq2885, weq2884, weq2883, weq2882, weq2881, weq2880, weq2879, weq2878, weq2877, weq2876, weq2875, weq2874, weq2873, weq2872, weq2871, weq2870, weq2869, weq2868, weq2867, weq2866, weq2865, weq2864, weq2863, weq2862, weq2861, weq2860, weq2859, weq2858, weq2857, weq2856, weq2855, weq2854, weq2853, weq2852, weq2851, weq2850, weq2849, weq2848, weq2847, weq2846, weq2845, weq2844, weq2843, weq2842, weq2841, weq2840, weq2839, weq2838, weq2837, weq2836, weq2835, weq2834, weq2833, weq2832, weq2831, weq2830, weq2829, weq2828, weq2827, weq2826, weq2825, weq2824, weq2823, weq2822, weq2821, weq2820, weq2819, weq2818, weq2817, weq2816, weq2815, weq2814, weq2813, weq2812, weq2811, weq2810, weq2809, weq2808, weq2807, weq2806, weq2805, weq2804, weq2803, weq2802, weq2801, weq2800, weq2799, weq2798, weq2797, weq2796, weq2795, weq2794, weq2793, weq2792, weq2791, weq2790, weq2789, weq2788, weq2787, weq2786, weq2785, weq2784, weq2783, weq2782, weq2781, weq2780, weq2779, weq2778, weq2777, weq2776, weq2775, weq2774, weq2773, weq2772, weq2771, weq2770, weq2769, weq2768, weq2767, weq2766, weq2765, weq2764, weq2763, weq2762, weq2761, weq2760, weq2759, weq2758, weq2757, weq2756, weq2755, weq2754, weq2753, weq2752, weq2751, weq2750, weq2749, weq2748, weq2747, weq2746, weq2745, weq2744, weq2743, weq2742, weq2741, weq2740, weq2739, weq2738, weq2737, weq2736, weq2735, weq2734, weq2733, weq2732, weq2731, weq2730, weq2729, weq2728, weq2727, weq2726, weq2725, weq2724, weq2723, weq2722, weq2721, weq2720, weq2719, weq2718, weq2717, weq2716, weq2715, weq2714, weq2713, weq2712, weq2711, weq2710, weq2709, weq2708, weq2707, weq2706, weq2705, weq2704, weq2703, weq2702, weq2701, weq2700, weq2699, weq2698, weq2697, weq2696, weq2695, weq2694, weq2693, weq2692, weq2691, weq2690, weq2689, weq2688, weq2687, weq2686, weq2685, weq2684, weq2683, weq2682, weq2681, weq2680, weq2679, weq2678, weq2677, weq2676, weq2675, weq2674, weq2673, weq2672, weq2671, weq2670, weq2669, weq2668, weq2667, weq2666, weq2665, weq2664, weq2663, weq2662, weq2661, weq2660, weq2659, weq2658, weq2657, weq2656, weq2655, weq2654, weq2653, weq2652, weq2651, weq2650, weq2649, weq2648, weq2647, weq2646, weq2645, weq2644, weq2643, weq2642, weq2641, weq2640, weq2639, weq2638, weq2637, weq2636, weq2635, weq2634, weq2633, weq2632, weq2631, weq2630, weq2629, weq2628, weq2627, weq2626, weq2625, weq2624, weq2623, weq2622, weq2621, weq2620, weq2619, weq2618, weq2617, weq2616, weq2615, weq2614, weq2613, weq2612, weq2611, weq2610, weq2609, weq2608, weq2607, weq2606, weq2605, weq2604, weq2603, weq2602, weq2601, weq2600, weq2599, weq2598, weq2597, weq2596, weq2595, weq2594, weq2593, weq2592, weq2591, weq2590, weq2589, weq2588, weq2587, weq2586, weq2585, weq2584, weq2583, weq2582, weq2581, weq2580, weq2579, weq2578, weq2577, weq2576, weq2575, weq2574, weq2573, weq2572, weq2571, weq2570, weq2569, weq2568, weq2567, weq2566, weq2565, weq2564, weq2563, weq2562, weq2561, weq2560, weq2559, weq2558, weq2557, weq2556, weq2555, weq2554, weq2553, weq2552, weq2551, weq2550, weq2549, weq2548, weq2547, weq2546, weq2545, weq2544, weq2543, weq2542, weq2541, weq2540, weq2539, weq2538, weq2537, weq2536, weq2535, weq2534, weq2533, weq2532, weq2531, weq2530, weq2529, weq2528, weq2527, weq2526, weq2525, weq2524, weq2523, weq2522, weq2521, weq2520, weq2519, weq2518, weq2517, weq2516, weq2515, weq2514, weq2513, weq2512, weq2511, weq2510, weq2509, weq2508, weq2507, weq2506, weq2505, weq2504, weq2503, weq2502, weq2501, weq2500, weq2499, weq2498, weq2497, weq2496, weq2495, weq2494, weq2493, weq2492, weq2491, weq2490, weq2489, weq2488, weq2487, weq2486, weq2485, weq2484, weq2483, weq2482, weq2481, weq2480, weq2479, weq2478, weq2477, weq2476, weq2475, weq2474, weq2473, weq2472, weq2471, weq2470, weq2469, weq2468, weq2467, weq2466, weq2465, weq2464, weq2463, weq2462, weq2461, weq2460, weq2459, weq2458, weq2457, weq2456, weq2455, weq2454, weq2453, weq2452, weq2451, weq2450, weq2449, weq2448, weq2447, weq2446, weq2445, weq2444, weq2443, weq2442, weq2441, weq2440, weq2439, weq2438, weq2437, weq2436, weq2435, weq2434, weq2433, weq2432, weq2431, weq2430, weq2429, weq2428, weq2427, weq2426, weq2425, weq2424, weq2423, weq2422, weq2421, weq2420, weq2419, weq2418, weq2417, weq2416, weq2415, weq2414, weq2413, weq2412, weq2411, weq2410, weq2409, weq2408, weq2407, weq2406, weq2405, weq2404, weq2403, weq2402, weq2401, weq2400, weq2399, weq2398, weq2397, weq2396, weq2395, weq2394, weq2393, weq2392, weq2391, weq2390, weq2389, weq2388, weq2387, weq2386, weq2385, weq2384, weq2383, weq2382, weq2381, weq2380, weq2379, weq2378, weq2377, weq2376, weq2375, weq2374, weq2373, weq2372, weq2371, weq2370, weq2369, weq2368, weq2367, weq2366, weq2365, weq2364, weq2363, weq2362, weq2361, weq2360, weq2359, weq2358, weq2357, weq2356, weq2355, weq2354, weq2353, weq2352, weq2351, weq2350, weq2349, weq2348, weq2347, weq2346, weq2345, weq2344, weq2343, weq2342, weq2341, weq2340, weq2339, weq2338, weq2337, weq2336, weq2335, weq2334, weq2333, weq2332, weq2331, weq2330, weq2329, weq2328, weq2327, weq2326, weq2325, weq2324, weq2323, weq2322, weq2321, weq2320, weq2319, weq2318, weq2317, weq2316, weq2315, weq2314, weq2313, weq2312, weq2311, weq2310, weq2309, weq2308, weq2307, weq2306, weq2305, weq2304, weq2303, weq2302, weq2301, weq2300, weq2299, weq2298, weq2297, weq2296, weq2295, weq2294, weq2293, weq2292, weq2291, weq2290, weq2289, weq2288, weq2287, weq2286, weq2285, weq2284, weq2283, weq2282, weq2281, weq2280, weq2279, weq2278, weq2277, weq2276, weq2275, weq2274, weq2273, weq2272, weq2271, weq2270, weq2269, weq2268, weq2267, weq2266, weq2265, weq2264, weq2263, weq2262, weq2261, weq2260, weq2259, weq2258, weq2257, weq2256, weq2255, weq2254, weq2253, weq2252, weq2251, weq2250, weq2249, weq2248, weq2247, weq2246, weq2245, weq2244, weq2243, weq2242, weq2241, weq2240, weq2239, weq2238, weq2237, weq2236, weq2235, weq2234, weq2233, weq2232, weq2231, weq2230, weq2229, weq2228, weq2227, weq2226, weq2225, weq2224, weq2223, weq2222, weq2221, weq2220, weq2219, weq2218, weq2217, weq2216, weq2215, weq2214, weq2213, weq2212, weq2211, weq2210, weq2209, weq2208, weq2207, weq2206, weq2205, weq2204, weq2203, weq2202, weq2201, weq2200, weq2199, weq2198, weq2197, weq2196, weq2195, weq2194, weq2193, weq2192, weq2191, weq2190, weq2189, weq2188, weq2187, weq2186, weq2185, weq2184, weq2183, weq2182, weq2181, weq2180, weq2179, weq2178, weq2177, weq2176, weq2175, weq2174, weq2173, weq2172, weq2171, weq2170, weq2169, weq2168, weq2167, weq2166, weq2165, weq2164, weq2163, weq2162, weq2161, weq2160, weq2159, weq2158, weq2157, weq2156, weq2155, weq2154, weq2153, weq2152, weq2151, weq2150, weq2149, weq2148, weq2147, weq2146, weq2145, weq2144, weq2143, weq2142, weq2141, weq2140, weq2139, weq2138, weq2137, weq2136, weq2135, weq2134, weq2133, weq2132, weq2131, weq2130, weq2129, weq2128, weq2127, weq2126, weq2125, weq2124, weq2123, weq2122, weq2121, weq2120, weq2119, weq2118, weq2117, weq2116, weq2115, weq2114, weq2113, weq2112, weq2111, weq2110, weq2109, weq2108, weq2107, weq2106, weq2105, weq2104, weq2103, weq2102, weq2101, weq2100, weq2099, weq2098, weq2097, weq2096, weq2095, weq2094, weq2093, weq2092, weq2091, weq2090, weq2089, weq2088, weq2087, weq2086, weq2085, weq2084, weq2083, weq2082, weq2081, weq2080, weq2079, weq2078, weq2077, weq2076, weq2075, weq2074, weq2073, weq2072, weq2071, weq2070, weq2069, weq2068, weq2067, weq2066, weq2065, weq2064, weq2063, weq2062, weq2061, weq2060, weq2059, weq2058, weq2057, weq2056, weq2055, weq2054, weq2053, weq2052, weq2051, weq2050, weq2049, weq2048, weq2047, weq2046, weq2045, weq2044, weq2043, weq2042, weq2041, weq2040, weq2039, weq2038, weq2037, weq2036, weq2035, weq2034, weq2033, weq2032, weq2031, weq2030, weq2029, weq2028, weq2027, weq2026, weq2025, weq2024, weq2023, weq2022, weq2021, weq2020, weq2019, weq2018, weq2017, weq2016, weq2015, weq2014, weq2013, weq2012, weq2011, weq2010, weq2009, weq2008, weq2007, weq2006, weq2005, weq2004, weq2003, weq2002, weq2001, weq2000, weq1999, weq1998, weq1997, weq1996, weq1995, weq1994, weq1993, weq1992, weq1991, weq1990, weq1989, weq1988, weq1987, weq1986, weq1985, weq1984, weq1983, weq1982, weq1981, weq1980, weq1979, weq1978, weq1977, weq1976, weq1975, weq1974, weq1973, weq1972, weq1971, weq1970, weq1969, weq1968, weq1967, weq1966, weq1965, weq1964, weq1963, weq1962, weq1961, weq1960, weq1959, weq1958, weq1957, weq1956, weq1955, weq1954, weq1953, weq1952, weq1951, weq1950, weq1949, weq1948, weq1947, weq1946, weq1945, weq1944, weq1943, weq1942, weq1941, weq1940, weq1939, weq1938, weq1937, weq1936, weq1935, weq1934, weq1933, weq1932, weq1931, weq1930, weq1929, weq1928, weq1927, weq1926, weq1925, weq1924, weq1923, weq1922, weq1921, weq1920, weq1919, weq1918, weq1917, weq1916, weq1915, weq1914, weq1913, weq1912, weq1911, weq1910, weq1909, weq1908, weq1907, weq1906, weq1905, weq1904, weq1903, weq1902, weq1901, weq1900, weq1899, weq1898, weq1897, weq1896, weq1895, weq1894, weq1893, weq1892, weq1891, weq1890, weq1889, weq1888, weq1887, weq1886, weq1885, weq1884, weq1883, weq1882, weq1881, weq1880, weq1879, weq1878, weq1877, weq1876, weq1875, weq1874, weq1873, weq1872, weq1871, weq1870, weq1869, weq1868, weq1867, weq1866, weq1865, weq1864, weq1863, weq1862, weq1861, weq1860, weq1859, weq1858, weq1857, weq1856, weq1855, weq1854, weq1853, weq1852, weq1851, weq1850, weq1849, weq1848, weq1847, weq1846, weq1845, weq1844, weq1843, weq1842, weq1841, weq1840, weq1839, weq1838, weq1837, weq1836, weq1835, weq1834, weq1833, weq1832, weq1831, weq1830, weq1829, weq1828, weq1827, weq1826, weq1825, weq1824, weq1823, weq1822, weq1821, weq1820, weq1819, weq1818, weq1817, weq1816, weq1815, weq1814, weq1813, weq1812, weq1811, weq1810, weq1809, weq1808, weq1807, weq1806, weq1805, weq1804, weq1803, weq1802, weq1801, weq1800, weq1799, weq1798, weq1797, weq1796, weq1795, weq1794, weq1793, weq1792, weq1791, weq1790, weq1789, weq1788, weq1787, weq1786, weq1785, weq1784, weq1783, weq1782, weq1781, weq1780, weq1779, weq1778, weq1777, weq1776, weq1775, weq1774, weq1773, weq1772, weq1771, weq1770, weq1769, weq1768, weq1767, weq1766, weq1765, weq1764, weq1763, weq1762, weq1761, weq1760, weq1759, weq1758, weq1757, weq1756, weq1755, weq1754, weq1753, weq1752, weq1751, weq1750, weq1749, weq1748, weq1747, weq1746, weq1745, weq1744, weq1743, weq1742, weq1741, weq1740, weq1739, weq1738, weq1737, weq1736, weq1735, weq1734, weq1733, weq1732, weq1731, weq1730, weq1729, weq1728, weq1727, weq1726, weq1725, weq1724, weq1723, weq1722, weq1721, weq1720, weq1719, weq1718, weq1717, weq1716, weq1715, weq1714, weq1713, weq1712, weq1711, weq1710, weq1709, weq1708, weq1707, weq1706, weq1705, weq1704, weq1703, weq1702, weq1701, weq1700, weq1699, weq1698, weq1697, weq1696, weq1695, weq1694, weq1693, weq1692, weq1691, weq1690, weq1689, weq1688, weq1687, weq1686, weq1685, weq1684, weq1683, weq1682, weq1681, weq1680, weq1679, weq1678, weq1677, weq1676, weq1675, weq1674, weq1673, weq1672, weq1671, weq1670, weq1669, weq1668, weq1667, weq1666, weq1665, weq1664, weq1663, weq1662, weq1661, weq1660, weq1659, weq1658, weq1657, weq1656, weq1655, weq1654, weq1653, weq1652, weq1651, weq1650, weq1649, weq1648, weq1647, weq1646, weq1645, weq1644, weq1643, weq1642, weq1641, weq1640, weq1639, weq1638, weq1637, weq1636, weq1635, weq1634, weq1633, weq1632, weq1631, weq1630, weq1629, weq1628, weq1627, weq1626, weq1625, weq1624, weq1623, weq1622, weq1621, weq1620, weq1619, weq1618, weq1617, weq1616, weq1615, weq1614, weq1613, weq1612, weq1611, weq1610, weq1609, weq1608, weq1607, weq1606, weq1605, weq1604, weq1603, weq1602, weq1601, weq1600, weq1599, weq1598, weq1597, weq1596, weq1595, weq1594, weq1593, weq1592, weq1591, weq1590, weq1589, weq1588, weq1587, weq1586, weq1585, weq1584, weq1583, weq1582, weq1581, weq1580, weq1579, weq1578, weq1577, weq1576, weq1575, weq1574, weq1573, weq1572, weq1571, weq1570, weq1569, weq1568, weq1567, weq1566, weq1565, weq1564, weq1563, weq1562, weq1561, weq1560, weq1559, weq1558, weq1557, weq1556, weq1555, weq1554, weq1553, weq1552, weq1551, weq1550, weq1549, weq1548, weq1547, weq1546, weq1545, weq1544, weq1543, weq1542, weq1541, weq1540, weq1539, weq1538, weq1537, weq1536, weq1535, weq1534, weq1533, weq1532, weq1531, weq1530, weq1529, weq1528, weq1527, weq1526, weq1525, weq1524, weq1523, weq1522, weq1521, weq1520, weq1519, weq1518, weq1517, weq1516, weq1515, weq1514, weq1513, weq1512, weq1511, weq1510, weq1509, weq1508, weq1507, weq1506, weq1505, weq1504, weq1503, weq1502, weq1501, weq1500, weq1499, weq1498, weq1497, weq1496, weq1495, weq1494, weq1493, weq1492, weq1491, weq1490, weq1489, weq1488, weq1487, weq1486, weq1485, weq1484, weq1483, weq1482, weq1481, weq1480, weq1479, weq1478, weq1477, weq1476, weq1475, weq1474, weq1473, weq1472, weq1471, weq1470, weq1469, weq1468, weq1467, weq1466, weq1465, weq1464, weq1463, weq1462, weq1461, weq1460, weq1459, weq1458, weq1457, weq1456, weq1455, weq1454, weq1453, weq1452, weq1451, weq1450, weq1449, weq1448, weq1447, weq1446, weq1445, weq1444, weq1443, weq1442, weq1441, weq1440, weq1439, weq1438, weq1437, weq1436, weq1435, weq1434, weq1433, weq1432, weq1431, weq1430, weq1429, weq1428, weq1427, weq1426, weq1425, weq1424, weq1423, weq1422, weq1421, weq1420, weq1419, weq1418, weq1417, weq1416, weq1415, weq1414, weq1413, weq1412, weq1411, weq1410, weq1409, weq1408, weq1407, weq1406, weq1405, weq1404, weq1403, weq1402, weq1401, weq1400, weq1399, weq1398, weq1397, weq1396, weq1395, weq1394, weq1393, weq1392, weq1391, weq1390, weq1389, weq1388, weq1387, weq1386, weq1385, weq1384, weq1383, weq1382, weq1381, weq1380, weq1379, weq1378, weq1377, weq1376, weq1375, weq1374, weq1373, weq1372, weq1371, weq1370, weq1369, weq1368, weq1367, weq1366, weq1365, weq1364, weq1363, weq1362, weq1361, weq1360, weq1359, weq1358, weq1357, weq1356, weq1355, weq1354, weq1353, weq1352, weq1351, weq1350, weq1349, weq1348, weq1347, weq1346, weq1345, weq1344, weq1343, weq1342, weq1341, weq1340, weq1339, weq1338, weq1337, weq1336, weq1335, weq1334, weq1333, weq1332, weq1331, weq1330, weq1329, weq1328, weq1327, weq1326, weq1325, weq1324, weq1323, weq1322, weq1321, weq1320, weq1319, weq1318, weq1317, weq1316, weq1315, weq1314, weq1313, weq1312, weq1311, weq1310, weq1309, weq1308, weq1307, weq1306, weq1305, weq1304, weq1303, weq1302, weq1301, weq1300, weq1299, weq1298, weq1297, weq1296, weq1295, weq1294, weq1293, weq1292, weq1291, weq1290, weq1289, weq1288, weq1287, weq1286, weq1285, weq1284, weq1283, weq1282, weq1281, weq1280, weq1279, weq1278, weq1277, weq1276, weq1275, weq1274, weq1273, weq1272, weq1271, weq1270, weq1269, weq1268, weq1267, weq1266, weq1265, weq1264, weq1263, weq1262, weq1261, weq1260, weq1259, weq1258, weq1257, weq1256, weq1255, weq1254, weq1253, weq1252, weq1251, weq1250, weq1249, weq1248, weq1247, weq1246, weq1245, weq1244, weq1243, weq1242, weq1241, weq1240, weq1239, weq1238, weq1237, weq1236, weq1235, weq1234, weq1233, weq1232, weq1231, weq1230, weq1229, weq1228, weq1227, weq1226, weq1225, weq1224, weq1223, weq1222, weq1221, weq1220, weq1219, weq1218, weq1217, weq1216, weq1215, weq1214, weq1213, weq1212, weq1211, weq1210, weq1209, weq1208, weq1207, weq1206, weq1205, weq1204, weq1203, weq1202, weq1201, weq1200, weq1199, weq1198, weq1197, weq1196, weq1195, weq1194, weq1193, weq1192, weq1191, weq1190, weq1189, weq1188, weq1187, weq1186, weq1185, weq1184, weq1183, weq1182, weq1181, weq1180, weq1179, weq1178, weq1177, weq1176, weq1175, weq1174, weq1173, weq1172, weq1171, weq1170, weq1169, weq1168, weq1167, weq1166, weq1165, weq1164, weq1163, weq1162, weq1161, weq1160, weq1159, weq1158, weq1157, weq1156, weq1155, weq1154, weq1153, weq1152, weq1151, weq1150, weq1149, weq1148, weq1147, weq1146, weq1145, weq1144, weq1143, weq1142, weq1141, weq1140, weq1139, weq1138, weq1137, weq1136, weq1135, weq1134, weq1133, weq1132, weq1131, weq1130, weq1129, weq1128, weq1127, weq1126, weq1125, weq1124, weq1123, weq1122, weq1121, weq1120, weq1119, weq1118, weq1117, weq1116, weq1115, weq1114, weq1113, weq1112, weq1111, weq1110, weq1109, weq1108, weq1107, weq1106, weq1105, weq1104, weq1103, weq1102, weq1101, weq1100, weq1099, weq1098, weq1097, weq1096, weq1095, weq1094, weq1093, weq1092, weq1091, weq1090, weq1089, weq1088, weq1087, weq1086, weq1085, weq1084, weq1083, weq1082, weq1081, weq1080, weq1079, weq1078, weq1077, weq1076, weq1075, weq1074, weq1073, weq1072, weq1071, weq1070, weq1069, weq1068, weq1067, weq1066, weq1065, weq1064, weq1063, weq1062, weq1061, weq1060, weq1059, weq1058, weq1057, weq1056, weq1055, weq1054, weq1053, weq1052, weq1051, weq1050, weq1049, weq1048, weq1047, weq1046, weq1045, weq1044, weq1043, weq1042, weq1041, weq1040, weq1039, weq1038, weq1037, weq1036, weq1035, weq1034, weq1033, weq1032, weq1031, weq1030, weq1029, weq1028, weq1027, weq1026, weq1025, weq1024, weq1023, weq1022, weq1021, weq1020, weq1019, weq1018, weq1017, weq1016, weq1015, weq1014, weq1013, weq1012, weq1011, weq1010, weq1009, weq1008, weq1007, weq1006, weq1005, weq1004, weq1003, weq1002, weq1001, weq1000, weq999, weq998, weq997, weq996, weq995, weq994, weq993, weq992, weq991, weq990, weq989, weq988, weq987, weq986, weq985, weq984, weq983, weq982, weq981, weq980, weq979, weq978, weq977, weq976, weq975, weq974, weq973, weq972, weq971, weq970, weq969, weq968, weq967, weq966, weq965, weq964, weq963, weq962, weq961, weq960, weq959, weq958, weq957, weq956, weq955, weq954, weq953, weq952, weq951, weq950, weq949, weq948, weq947, weq946, weq945, weq944, weq943, weq942, weq941, weq940, weq939, weq938, weq937, weq936, weq935, weq934, weq933, weq932, weq931, weq930, weq929, weq928, weq927, weq926, weq925, weq924, weq923, weq922, weq921, weq920, weq919, weq918, weq917, weq916, weq915, weq914, weq913, weq912, weq911, weq910, weq909, weq908, weq907, weq906, weq905, weq904, weq903, weq902, weq901, weq900, weq899, weq898, weq897, weq896, weq895, weq894, weq893, weq892, weq891, weq890, weq889, weq888, weq887, weq886, weq885, weq884, weq883, weq882, weq881, weq880, weq879, weq878, weq877, weq876, weq875, weq874, weq873, weq872, weq871, weq870, weq869, weq868, weq867, weq866, weq865, weq864, weq863, weq862, weq861, weq860, weq859, weq858, weq857, weq856, weq855, weq854, weq853, weq852, weq851, weq850, weq849, weq848, weq847, weq846, weq845, weq844, weq843, weq842, weq841, weq840, weq839, weq838, weq837, weq836, weq835, weq834, weq833, weq832, weq831, weq830, weq829, weq828, weq827, weq826, weq825, weq824, weq823, weq822, weq821, weq820, weq819, weq818, weq817, weq816, weq815, weq814, weq813, weq812, weq811, weq810, weq809, weq808, weq807, weq806, weq805, weq804, weq803, weq802, weq801, weq800, weq799, weq798, weq797, weq796, weq795, weq794, weq793, weq792, weq791, weq790, weq789, weq788, weq787, weq786, weq785, weq784, weq783, weq782, weq781, weq780, weq779, weq778, weq777, weq776, weq775, weq774, weq773, weq772, weq771, weq770, weq769, weq768, weq767, weq766, weq765, weq764, weq763, weq762, weq761, weq760, weq759, weq758, weq757, weq756, weq755, weq754, weq753, weq752, weq751, weq750, weq749, weq748, weq747, weq746, weq745, weq744, weq743, weq742, weq741, weq740, weq739, weq738, weq737, weq736, weq735, weq734, weq733, weq732, weq731, weq730, weq729, weq728, weq727, weq726, weq725, weq724, weq723, weq722, weq721, weq720, weq719, weq718, weq717, weq716, weq715, weq714, weq713, weq712, weq711, weq710, weq709, weq708, weq707, weq706, weq705, weq704, weq703, weq702, weq701, weq700, weq699, weq698, weq697, weq696, weq695, weq694, weq693, weq692, weq691, weq690, weq689, weq688, weq687, weq686, weq685, weq684, weq683, weq682, weq681, weq680, weq679, weq678, weq677, weq676, weq675, weq674, weq673, weq672, weq671, weq670, weq669, weq668, weq667, weq666, weq665, weq664, weq663, weq662, weq661, weq660, weq659, weq658, weq657, weq656, weq655, weq654, weq653, weq652, weq651, weq650, weq649, weq648, weq647, weq646, weq645, weq644, weq643, weq642, weq641, weq640, weq639, weq638, weq637, weq636, weq635, weq634, weq633, weq632, weq631, weq630, weq629, weq628, weq627, weq626, weq625, weq624, weq623, weq622, weq621, weq620, weq619, weq618, weq617, weq616, weq615, weq614, weq613, weq612, weq611, weq610, weq609, weq608, weq607, weq606, weq605, weq604, weq603, weq602, weq601, weq600, weq599, weq598, weq597, weq596, weq595, weq594, weq593, weq592, weq591, weq590, weq589, weq588, weq587, weq586, weq585, weq584, weq583, weq582, weq581, weq580, weq579, weq578, weq577, weq576, weq575, weq574, weq573, weq572, weq571, weq570, weq569, weq568, weq567, weq566, weq565, weq564, weq563, weq562, weq561, weq560, weq559, weq558, weq557, weq556, weq555, weq554, weq553, weq552, weq551, weq550, weq549, weq548, weq547, weq546, weq545, weq544, weq543, weq542, weq541, weq540, weq539, weq538, weq537, weq536, weq535, weq534, weq533, weq532, weq531, weq530, weq529, weq528, weq527, weq526, weq525, weq524, weq523, weq522, weq521, weq520, weq519, weq518, weq517, weq516, weq515, weq514, weq513, weq512, weq511, weq510, weq509, weq508, weq507, weq506, weq505, weq504, weq503, weq502, weq501, weq500, weq499, weq498, weq497, weq496, weq495, weq494, weq493, weq492, weq491, weq490, weq489, weq488, weq487, weq486, weq485, weq484, weq483, weq482, weq481, weq480, weq479, weq478, weq477, weq476, weq475, weq474, weq473, weq472, weq471, weq470, weq469, weq468, weq467, weq466, weq465, weq464, weq463, weq462, weq461, weq460, weq459, weq458, weq457, weq456, weq455, weq454, weq453, weq452, weq451, weq450, weq449, weq448, weq447, weq446, weq445, weq444, weq443, weq442, weq441, weq440, weq439, weq438, weq437, weq436, weq435, weq434, weq433, weq432, weq431, weq430, weq429, weq428, weq427, weq426, weq425, weq424, weq423, weq422, weq421, weq420, weq419, weq418, weq417, weq416, weq415, weq414, weq413, weq412, weq411, weq410, weq409, weq408, weq407, weq406, weq405, weq404, weq403, weq402, weq401, weq400, weq399, weq398, weq397, weq396, weq395, weq394, weq393, weq392, weq391, weq390, weq389, weq388, weq387, weq386, weq385, weq384, weq383, weq382, weq381, weq380, weq379, weq378, weq377, weq376, weq375, weq374, weq373, weq372, weq371, weq370, weq369, weq368, weq367, weq366, weq365, weq364, weq363, weq362, weq361, weq360, weq359, weq358, weq357, weq356, weq355, weq354, weq353, weq352, weq351, weq350, weq349, weq348, weq347, weq346, weq345, weq344, weq343, weq342, weq341, weq340, weq339, weq338, weq337, weq336, weq335, weq334, weq333, weq332, weq331, weq330, weq329, weq328, weq327, weq326, weq325, weq324, weq323, weq322, weq321, weq320, weq319, weq318, weq317, weq316, weq315, weq314, weq313, weq312, weq311, weq310, weq309, weq308, weq307, weq306, weq305, weq304, weq303, weq302, weq301, weq300, weq299, weq298, weq297, weq296, weq295, weq294, weq293, weq292, weq291, weq290, weq289, weq288, weq287, weq286, weq285, weq284, weq283, weq282, weq281, weq280, weq279, weq278, weq277, weq276, weq275, weq274, weq273, weq272, weq271, weq270, weq269, weq268, weq267, weq266, weq265, weq264, weq263, weq262, weq261, weq260, weq259, weq258, weq257, weq256, weq255, weq254, weq253, weq252, weq251, weq250, weq249, weq248, weq247, weq246, weq245, weq244, weq243, weq242, weq241, weq240, weq239, weq238, weq237, weq236, weq235, weq234, weq233, weq232, weq231, weq230, weq229, weq228, weq227, weq226, weq225, weq224, weq223, weq222, weq221, weq220, weq219, weq218, weq217, weq216, weq215, weq214, weq213, weq212, weq211, weq210, weq209, weq208, weq207, weq206, weq205, weq204, weq203, weq202, weq201, weq200, weq199, weq198, weq197, weq196, weq195, weq194, weq193, weq192, weq191, weq190, weq189, weq188, weq187, weq186, weq185, weq184, weq183, weq182, weq181, weq180, weq179, weq178, weq177, weq176, weq175, weq174, weq173, weq172, weq171, weq170, weq169, weq168, weq167, weq166, weq165, weq164, weq163, weq162, weq161, weq160, weq159, weq158, weq157, weq156, weq155, weq154, weq153, weq152, weq151, weq150, weq149, weq148, weq147, weq146, weq145, weq144, weq143, weq142, weq141, weq140, weq139, weq138, weq137, weq136, weq135, weq134, weq133, weq132, weq131, weq130, weq129, weq128, weq127, weq126, weq125, weq124, weq123, weq122, weq121, weq120, weq119, weq118, weq117, weq116, weq115, weq114, weq113, weq112, weq111, weq110, weq109, weq108, weq107, weq106, weq105, weq104, weq103, weq102, weq101, weq100, weq99, weq98, weq97, weq96, weq95, weq94, weq93, weq92, weq91, weq90, weq89, weq88, weq87, weq86, weq85, weq84, weq83, weq82, weq81, weq80, weq79, weq78, weq77, weq76, weq75, weq74, weq73, weq72, weq71, weq70, weq69, weq68, weq67, weq66, weq65, weq64, weq63, weq62, weq61, weq60, weq59, weq58, weq57, weq56, weq55, weq54, weq53, weq52, weq51, weq50, weq49, weq48, weq47, weq46, weq45, weq44, weq43, weq42, weq41, weq40, weq39, weq38, weq37, weq36, weq35, weq34, weq33, weq32, weq31, weq30, weq29, weq28, weq27, weq26, weq25, weq24, weq23, weq22, weq21, weq20, weq19, weq18, weq17, weq16, weq15, weq14, weq13, weq12, weq11, weq10, weq9, weq8, weq7, weq6, weq5, weq4, weq3, weq2, weq1, weq0};

    wire [32767:0] data_concat;
    assign data_concat = {wire4095, wire4094, wire4093, wire4092, wire4091, wire4090, wire4089, wire4088, wire4087, wire4086, wire4085, wire4084, wire4083, wire4082, wire4081, wire4080, wire4079, wire4078, wire4077, wire4076, wire4075, wire4074, wire4073, wire4072, wire4071, wire4070, wire4069, wire4068, wire4067, wire4066, wire4065, wire4064, wire4063, wire4062, wire4061, wire4060, wire4059, wire4058, wire4057, wire4056, wire4055, wire4054, wire4053, wire4052, wire4051, wire4050, wire4049, wire4048, wire4047, wire4046, wire4045, wire4044, wire4043, wire4042, wire4041, wire4040, wire4039, wire4038, wire4037, wire4036, wire4035, wire4034, wire4033, wire4032, wire4031, wire4030, wire4029, wire4028, wire4027, wire4026, wire4025, wire4024, wire4023, wire4022, wire4021, wire4020, wire4019, wire4018, wire4017, wire4016, wire4015, wire4014, wire4013, wire4012, wire4011, wire4010, wire4009, wire4008, wire4007, wire4006, wire4005, wire4004, wire4003, wire4002, wire4001, wire4000, wire3999, wire3998, wire3997, wire3996, wire3995, wire3994, wire3993, wire3992, wire3991, wire3990, wire3989, wire3988, wire3987, wire3986, wire3985, wire3984, wire3983, wire3982, wire3981, wire3980, wire3979, wire3978, wire3977, wire3976, wire3975, wire3974, wire3973, wire3972, wire3971, wire3970, wire3969, wire3968, wire3967, wire3966, wire3965, wire3964, wire3963, wire3962, wire3961, wire3960, wire3959, wire3958, wire3957, wire3956, wire3955, wire3954, wire3953, wire3952, wire3951, wire3950, wire3949, wire3948, wire3947, wire3946, wire3945, wire3944, wire3943, wire3942, wire3941, wire3940, wire3939, wire3938, wire3937, wire3936, wire3935, wire3934, wire3933, wire3932, wire3931, wire3930, wire3929, wire3928, wire3927, wire3926, wire3925, wire3924, wire3923, wire3922, wire3921, wire3920, wire3919, wire3918, wire3917, wire3916, wire3915, wire3914, wire3913, wire3912, wire3911, wire3910, wire3909, wire3908, wire3907, wire3906, wire3905, wire3904, wire3903, wire3902, wire3901, wire3900, wire3899, wire3898, wire3897, wire3896, wire3895, wire3894, wire3893, wire3892, wire3891, wire3890, wire3889, wire3888, wire3887, wire3886, wire3885, wire3884, wire3883, wire3882, wire3881, wire3880, wire3879, wire3878, wire3877, wire3876, wire3875, wire3874, wire3873, wire3872, wire3871, wire3870, wire3869, wire3868, wire3867, wire3866, wire3865, wire3864, wire3863, wire3862, wire3861, wire3860, wire3859, wire3858, wire3857, wire3856, wire3855, wire3854, wire3853, wire3852, wire3851, wire3850, wire3849, wire3848, wire3847, wire3846, wire3845, wire3844, wire3843, wire3842, wire3841, wire3840, wire3839, wire3838, wire3837, wire3836, wire3835, wire3834, wire3833, wire3832, wire3831, wire3830, wire3829, wire3828, wire3827, wire3826, wire3825, wire3824, wire3823, wire3822, wire3821, wire3820, wire3819, wire3818, wire3817, wire3816, wire3815, wire3814, wire3813, wire3812, wire3811, wire3810, wire3809, wire3808, wire3807, wire3806, wire3805, wire3804, wire3803, wire3802, wire3801, wire3800, wire3799, wire3798, wire3797, wire3796, wire3795, wire3794, wire3793, wire3792, wire3791, wire3790, wire3789, wire3788, wire3787, wire3786, wire3785, wire3784, wire3783, wire3782, wire3781, wire3780, wire3779, wire3778, wire3777, wire3776, wire3775, wire3774, wire3773, wire3772, wire3771, wire3770, wire3769, wire3768, wire3767, wire3766, wire3765, wire3764, wire3763, wire3762, wire3761, wire3760, wire3759, wire3758, wire3757, wire3756, wire3755, wire3754, wire3753, wire3752, wire3751, wire3750, wire3749, wire3748, wire3747, wire3746, wire3745, wire3744, wire3743, wire3742, wire3741, wire3740, wire3739, wire3738, wire3737, wire3736, wire3735, wire3734, wire3733, wire3732, wire3731, wire3730, wire3729, wire3728, wire3727, wire3726, wire3725, wire3724, wire3723, wire3722, wire3721, wire3720, wire3719, wire3718, wire3717, wire3716, wire3715, wire3714, wire3713, wire3712, wire3711, wire3710, wire3709, wire3708, wire3707, wire3706, wire3705, wire3704, wire3703, wire3702, wire3701, wire3700, wire3699, wire3698, wire3697, wire3696, wire3695, wire3694, wire3693, wire3692, wire3691, wire3690, wire3689, wire3688, wire3687, wire3686, wire3685, wire3684, wire3683, wire3682, wire3681, wire3680, wire3679, wire3678, wire3677, wire3676, wire3675, wire3674, wire3673, wire3672, wire3671, wire3670, wire3669, wire3668, wire3667, wire3666, wire3665, wire3664, wire3663, wire3662, wire3661, wire3660, wire3659, wire3658, wire3657, wire3656, wire3655, wire3654, wire3653, wire3652, wire3651, wire3650, wire3649, wire3648, wire3647, wire3646, wire3645, wire3644, wire3643, wire3642, wire3641, wire3640, wire3639, wire3638, wire3637, wire3636, wire3635, wire3634, wire3633, wire3632, wire3631, wire3630, wire3629, wire3628, wire3627, wire3626, wire3625, wire3624, wire3623, wire3622, wire3621, wire3620, wire3619, wire3618, wire3617, wire3616, wire3615, wire3614, wire3613, wire3612, wire3611, wire3610, wire3609, wire3608, wire3607, wire3606, wire3605, wire3604, wire3603, wire3602, wire3601, wire3600, wire3599, wire3598, wire3597, wire3596, wire3595, wire3594, wire3593, wire3592, wire3591, wire3590, wire3589, wire3588, wire3587, wire3586, wire3585, wire3584, wire3583, wire3582, wire3581, wire3580, wire3579, wire3578, wire3577, wire3576, wire3575, wire3574, wire3573, wire3572, wire3571, wire3570, wire3569, wire3568, wire3567, wire3566, wire3565, wire3564, wire3563, wire3562, wire3561, wire3560, wire3559, wire3558, wire3557, wire3556, wire3555, wire3554, wire3553, wire3552, wire3551, wire3550, wire3549, wire3548, wire3547, wire3546, wire3545, wire3544, wire3543, wire3542, wire3541, wire3540, wire3539, wire3538, wire3537, wire3536, wire3535, wire3534, wire3533, wire3532, wire3531, wire3530, wire3529, wire3528, wire3527, wire3526, wire3525, wire3524, wire3523, wire3522, wire3521, wire3520, wire3519, wire3518, wire3517, wire3516, wire3515, wire3514, wire3513, wire3512, wire3511, wire3510, wire3509, wire3508, wire3507, wire3506, wire3505, wire3504, wire3503, wire3502, wire3501, wire3500, wire3499, wire3498, wire3497, wire3496, wire3495, wire3494, wire3493, wire3492, wire3491, wire3490, wire3489, wire3488, wire3487, wire3486, wire3485, wire3484, wire3483, wire3482, wire3481, wire3480, wire3479, wire3478, wire3477, wire3476, wire3475, wire3474, wire3473, wire3472, wire3471, wire3470, wire3469, wire3468, wire3467, wire3466, wire3465, wire3464, wire3463, wire3462, wire3461, wire3460, wire3459, wire3458, wire3457, wire3456, wire3455, wire3454, wire3453, wire3452, wire3451, wire3450, wire3449, wire3448, wire3447, wire3446, wire3445, wire3444, wire3443, wire3442, wire3441, wire3440, wire3439, wire3438, wire3437, wire3436, wire3435, wire3434, wire3433, wire3432, wire3431, wire3430, wire3429, wire3428, wire3427, wire3426, wire3425, wire3424, wire3423, wire3422, wire3421, wire3420, wire3419, wire3418, wire3417, wire3416, wire3415, wire3414, wire3413, wire3412, wire3411, wire3410, wire3409, wire3408, wire3407, wire3406, wire3405, wire3404, wire3403, wire3402, wire3401, wire3400, wire3399, wire3398, wire3397, wire3396, wire3395, wire3394, wire3393, wire3392, wire3391, wire3390, wire3389, wire3388, wire3387, wire3386, wire3385, wire3384, wire3383, wire3382, wire3381, wire3380, wire3379, wire3378, wire3377, wire3376, wire3375, wire3374, wire3373, wire3372, wire3371, wire3370, wire3369, wire3368, wire3367, wire3366, wire3365, wire3364, wire3363, wire3362, wire3361, wire3360, wire3359, wire3358, wire3357, wire3356, wire3355, wire3354, wire3353, wire3352, wire3351, wire3350, wire3349, wire3348, wire3347, wire3346, wire3345, wire3344, wire3343, wire3342, wire3341, wire3340, wire3339, wire3338, wire3337, wire3336, wire3335, wire3334, wire3333, wire3332, wire3331, wire3330, wire3329, wire3328, wire3327, wire3326, wire3325, wire3324, wire3323, wire3322, wire3321, wire3320, wire3319, wire3318, wire3317, wire3316, wire3315, wire3314, wire3313, wire3312, wire3311, wire3310, wire3309, wire3308, wire3307, wire3306, wire3305, wire3304, wire3303, wire3302, wire3301, wire3300, wire3299, wire3298, wire3297, wire3296, wire3295, wire3294, wire3293, wire3292, wire3291, wire3290, wire3289, wire3288, wire3287, wire3286, wire3285, wire3284, wire3283, wire3282, wire3281, wire3280, wire3279, wire3278, wire3277, wire3276, wire3275, wire3274, wire3273, wire3272, wire3271, wire3270, wire3269, wire3268, wire3267, wire3266, wire3265, wire3264, wire3263, wire3262, wire3261, wire3260, wire3259, wire3258, wire3257, wire3256, wire3255, wire3254, wire3253, wire3252, wire3251, wire3250, wire3249, wire3248, wire3247, wire3246, wire3245, wire3244, wire3243, wire3242, wire3241, wire3240, wire3239, wire3238, wire3237, wire3236, wire3235, wire3234, wire3233, wire3232, wire3231, wire3230, wire3229, wire3228, wire3227, wire3226, wire3225, wire3224, wire3223, wire3222, wire3221, wire3220, wire3219, wire3218, wire3217, wire3216, wire3215, wire3214, wire3213, wire3212, wire3211, wire3210, wire3209, wire3208, wire3207, wire3206, wire3205, wire3204, wire3203, wire3202, wire3201, wire3200, wire3199, wire3198, wire3197, wire3196, wire3195, wire3194, wire3193, wire3192, wire3191, wire3190, wire3189, wire3188, wire3187, wire3186, wire3185, wire3184, wire3183, wire3182, wire3181, wire3180, wire3179, wire3178, wire3177, wire3176, wire3175, wire3174, wire3173, wire3172, wire3171, wire3170, wire3169, wire3168, wire3167, wire3166, wire3165, wire3164, wire3163, wire3162, wire3161, wire3160, wire3159, wire3158, wire3157, wire3156, wire3155, wire3154, wire3153, wire3152, wire3151, wire3150, wire3149, wire3148, wire3147, wire3146, wire3145, wire3144, wire3143, wire3142, wire3141, wire3140, wire3139, wire3138, wire3137, wire3136, wire3135, wire3134, wire3133, wire3132, wire3131, wire3130, wire3129, wire3128, wire3127, wire3126, wire3125, wire3124, wire3123, wire3122, wire3121, wire3120, wire3119, wire3118, wire3117, wire3116, wire3115, wire3114, wire3113, wire3112, wire3111, wire3110, wire3109, wire3108, wire3107, wire3106, wire3105, wire3104, wire3103, wire3102, wire3101, wire3100, wire3099, wire3098, wire3097, wire3096, wire3095, wire3094, wire3093, wire3092, wire3091, wire3090, wire3089, wire3088, wire3087, wire3086, wire3085, wire3084, wire3083, wire3082, wire3081, wire3080, wire3079, wire3078, wire3077, wire3076, wire3075, wire3074, wire3073, wire3072, wire3071, wire3070, wire3069, wire3068, wire3067, wire3066, wire3065, wire3064, wire3063, wire3062, wire3061, wire3060, wire3059, wire3058, wire3057, wire3056, wire3055, wire3054, wire3053, wire3052, wire3051, wire3050, wire3049, wire3048, wire3047, wire3046, wire3045, wire3044, wire3043, wire3042, wire3041, wire3040, wire3039, wire3038, wire3037, wire3036, wire3035, wire3034, wire3033, wire3032, wire3031, wire3030, wire3029, wire3028, wire3027, wire3026, wire3025, wire3024, wire3023, wire3022, wire3021, wire3020, wire3019, wire3018, wire3017, wire3016, wire3015, wire3014, wire3013, wire3012, wire3011, wire3010, wire3009, wire3008, wire3007, wire3006, wire3005, wire3004, wire3003, wire3002, wire3001, wire3000, wire2999, wire2998, wire2997, wire2996, wire2995, wire2994, wire2993, wire2992, wire2991, wire2990, wire2989, wire2988, wire2987, wire2986, wire2985, wire2984, wire2983, wire2982, wire2981, wire2980, wire2979, wire2978, wire2977, wire2976, wire2975, wire2974, wire2973, wire2972, wire2971, wire2970, wire2969, wire2968, wire2967, wire2966, wire2965, wire2964, wire2963, wire2962, wire2961, wire2960, wire2959, wire2958, wire2957, wire2956, wire2955, wire2954, wire2953, wire2952, wire2951, wire2950, wire2949, wire2948, wire2947, wire2946, wire2945, wire2944, wire2943, wire2942, wire2941, wire2940, wire2939, wire2938, wire2937, wire2936, wire2935, wire2934, wire2933, wire2932, wire2931, wire2930, wire2929, wire2928, wire2927, wire2926, wire2925, wire2924, wire2923, wire2922, wire2921, wire2920, wire2919, wire2918, wire2917, wire2916, wire2915, wire2914, wire2913, wire2912, wire2911, wire2910, wire2909, wire2908, wire2907, wire2906, wire2905, wire2904, wire2903, wire2902, wire2901, wire2900, wire2899, wire2898, wire2897, wire2896, wire2895, wire2894, wire2893, wire2892, wire2891, wire2890, wire2889, wire2888, wire2887, wire2886, wire2885, wire2884, wire2883, wire2882, wire2881, wire2880, wire2879, wire2878, wire2877, wire2876, wire2875, wire2874, wire2873, wire2872, wire2871, wire2870, wire2869, wire2868, wire2867, wire2866, wire2865, wire2864, wire2863, wire2862, wire2861, wire2860, wire2859, wire2858, wire2857, wire2856, wire2855, wire2854, wire2853, wire2852, wire2851, wire2850, wire2849, wire2848, wire2847, wire2846, wire2845, wire2844, wire2843, wire2842, wire2841, wire2840, wire2839, wire2838, wire2837, wire2836, wire2835, wire2834, wire2833, wire2832, wire2831, wire2830, wire2829, wire2828, wire2827, wire2826, wire2825, wire2824, wire2823, wire2822, wire2821, wire2820, wire2819, wire2818, wire2817, wire2816, wire2815, wire2814, wire2813, wire2812, wire2811, wire2810, wire2809, wire2808, wire2807, wire2806, wire2805, wire2804, wire2803, wire2802, wire2801, wire2800, wire2799, wire2798, wire2797, wire2796, wire2795, wire2794, wire2793, wire2792, wire2791, wire2790, wire2789, wire2788, wire2787, wire2786, wire2785, wire2784, wire2783, wire2782, wire2781, wire2780, wire2779, wire2778, wire2777, wire2776, wire2775, wire2774, wire2773, wire2772, wire2771, wire2770, wire2769, wire2768, wire2767, wire2766, wire2765, wire2764, wire2763, wire2762, wire2761, wire2760, wire2759, wire2758, wire2757, wire2756, wire2755, wire2754, wire2753, wire2752, wire2751, wire2750, wire2749, wire2748, wire2747, wire2746, wire2745, wire2744, wire2743, wire2742, wire2741, wire2740, wire2739, wire2738, wire2737, wire2736, wire2735, wire2734, wire2733, wire2732, wire2731, wire2730, wire2729, wire2728, wire2727, wire2726, wire2725, wire2724, wire2723, wire2722, wire2721, wire2720, wire2719, wire2718, wire2717, wire2716, wire2715, wire2714, wire2713, wire2712, wire2711, wire2710, wire2709, wire2708, wire2707, wire2706, wire2705, wire2704, wire2703, wire2702, wire2701, wire2700, wire2699, wire2698, wire2697, wire2696, wire2695, wire2694, wire2693, wire2692, wire2691, wire2690, wire2689, wire2688, wire2687, wire2686, wire2685, wire2684, wire2683, wire2682, wire2681, wire2680, wire2679, wire2678, wire2677, wire2676, wire2675, wire2674, wire2673, wire2672, wire2671, wire2670, wire2669, wire2668, wire2667, wire2666, wire2665, wire2664, wire2663, wire2662, wire2661, wire2660, wire2659, wire2658, wire2657, wire2656, wire2655, wire2654, wire2653, wire2652, wire2651, wire2650, wire2649, wire2648, wire2647, wire2646, wire2645, wire2644, wire2643, wire2642, wire2641, wire2640, wire2639, wire2638, wire2637, wire2636, wire2635, wire2634, wire2633, wire2632, wire2631, wire2630, wire2629, wire2628, wire2627, wire2626, wire2625, wire2624, wire2623, wire2622, wire2621, wire2620, wire2619, wire2618, wire2617, wire2616, wire2615, wire2614, wire2613, wire2612, wire2611, wire2610, wire2609, wire2608, wire2607, wire2606, wire2605, wire2604, wire2603, wire2602, wire2601, wire2600, wire2599, wire2598, wire2597, wire2596, wire2595, wire2594, wire2593, wire2592, wire2591, wire2590, wire2589, wire2588, wire2587, wire2586, wire2585, wire2584, wire2583, wire2582, wire2581, wire2580, wire2579, wire2578, wire2577, wire2576, wire2575, wire2574, wire2573, wire2572, wire2571, wire2570, wire2569, wire2568, wire2567, wire2566, wire2565, wire2564, wire2563, wire2562, wire2561, wire2560, wire2559, wire2558, wire2557, wire2556, wire2555, wire2554, wire2553, wire2552, wire2551, wire2550, wire2549, wire2548, wire2547, wire2546, wire2545, wire2544, wire2543, wire2542, wire2541, wire2540, wire2539, wire2538, wire2537, wire2536, wire2535, wire2534, wire2533, wire2532, wire2531, wire2530, wire2529, wire2528, wire2527, wire2526, wire2525, wire2524, wire2523, wire2522, wire2521, wire2520, wire2519, wire2518, wire2517, wire2516, wire2515, wire2514, wire2513, wire2512, wire2511, wire2510, wire2509, wire2508, wire2507, wire2506, wire2505, wire2504, wire2503, wire2502, wire2501, wire2500, wire2499, wire2498, wire2497, wire2496, wire2495, wire2494, wire2493, wire2492, wire2491, wire2490, wire2489, wire2488, wire2487, wire2486, wire2485, wire2484, wire2483, wire2482, wire2481, wire2480, wire2479, wire2478, wire2477, wire2476, wire2475, wire2474, wire2473, wire2472, wire2471, wire2470, wire2469, wire2468, wire2467, wire2466, wire2465, wire2464, wire2463, wire2462, wire2461, wire2460, wire2459, wire2458, wire2457, wire2456, wire2455, wire2454, wire2453, wire2452, wire2451, wire2450, wire2449, wire2448, wire2447, wire2446, wire2445, wire2444, wire2443, wire2442, wire2441, wire2440, wire2439, wire2438, wire2437, wire2436, wire2435, wire2434, wire2433, wire2432, wire2431, wire2430, wire2429, wire2428, wire2427, wire2426, wire2425, wire2424, wire2423, wire2422, wire2421, wire2420, wire2419, wire2418, wire2417, wire2416, wire2415, wire2414, wire2413, wire2412, wire2411, wire2410, wire2409, wire2408, wire2407, wire2406, wire2405, wire2404, wire2403, wire2402, wire2401, wire2400, wire2399, wire2398, wire2397, wire2396, wire2395, wire2394, wire2393, wire2392, wire2391, wire2390, wire2389, wire2388, wire2387, wire2386, wire2385, wire2384, wire2383, wire2382, wire2381, wire2380, wire2379, wire2378, wire2377, wire2376, wire2375, wire2374, wire2373, wire2372, wire2371, wire2370, wire2369, wire2368, wire2367, wire2366, wire2365, wire2364, wire2363, wire2362, wire2361, wire2360, wire2359, wire2358, wire2357, wire2356, wire2355, wire2354, wire2353, wire2352, wire2351, wire2350, wire2349, wire2348, wire2347, wire2346, wire2345, wire2344, wire2343, wire2342, wire2341, wire2340, wire2339, wire2338, wire2337, wire2336, wire2335, wire2334, wire2333, wire2332, wire2331, wire2330, wire2329, wire2328, wire2327, wire2326, wire2325, wire2324, wire2323, wire2322, wire2321, wire2320, wire2319, wire2318, wire2317, wire2316, wire2315, wire2314, wire2313, wire2312, wire2311, wire2310, wire2309, wire2308, wire2307, wire2306, wire2305, wire2304, wire2303, wire2302, wire2301, wire2300, wire2299, wire2298, wire2297, wire2296, wire2295, wire2294, wire2293, wire2292, wire2291, wire2290, wire2289, wire2288, wire2287, wire2286, wire2285, wire2284, wire2283, wire2282, wire2281, wire2280, wire2279, wire2278, wire2277, wire2276, wire2275, wire2274, wire2273, wire2272, wire2271, wire2270, wire2269, wire2268, wire2267, wire2266, wire2265, wire2264, wire2263, wire2262, wire2261, wire2260, wire2259, wire2258, wire2257, wire2256, wire2255, wire2254, wire2253, wire2252, wire2251, wire2250, wire2249, wire2248, wire2247, wire2246, wire2245, wire2244, wire2243, wire2242, wire2241, wire2240, wire2239, wire2238, wire2237, wire2236, wire2235, wire2234, wire2233, wire2232, wire2231, wire2230, wire2229, wire2228, wire2227, wire2226, wire2225, wire2224, wire2223, wire2222, wire2221, wire2220, wire2219, wire2218, wire2217, wire2216, wire2215, wire2214, wire2213, wire2212, wire2211, wire2210, wire2209, wire2208, wire2207, wire2206, wire2205, wire2204, wire2203, wire2202, wire2201, wire2200, wire2199, wire2198, wire2197, wire2196, wire2195, wire2194, wire2193, wire2192, wire2191, wire2190, wire2189, wire2188, wire2187, wire2186, wire2185, wire2184, wire2183, wire2182, wire2181, wire2180, wire2179, wire2178, wire2177, wire2176, wire2175, wire2174, wire2173, wire2172, wire2171, wire2170, wire2169, wire2168, wire2167, wire2166, wire2165, wire2164, wire2163, wire2162, wire2161, wire2160, wire2159, wire2158, wire2157, wire2156, wire2155, wire2154, wire2153, wire2152, wire2151, wire2150, wire2149, wire2148, wire2147, wire2146, wire2145, wire2144, wire2143, wire2142, wire2141, wire2140, wire2139, wire2138, wire2137, wire2136, wire2135, wire2134, wire2133, wire2132, wire2131, wire2130, wire2129, wire2128, wire2127, wire2126, wire2125, wire2124, wire2123, wire2122, wire2121, wire2120, wire2119, wire2118, wire2117, wire2116, wire2115, wire2114, wire2113, wire2112, wire2111, wire2110, wire2109, wire2108, wire2107, wire2106, wire2105, wire2104, wire2103, wire2102, wire2101, wire2100, wire2099, wire2098, wire2097, wire2096, wire2095, wire2094, wire2093, wire2092, wire2091, wire2090, wire2089, wire2088, wire2087, wire2086, wire2085, wire2084, wire2083, wire2082, wire2081, wire2080, wire2079, wire2078, wire2077, wire2076, wire2075, wire2074, wire2073, wire2072, wire2071, wire2070, wire2069, wire2068, wire2067, wire2066, wire2065, wire2064, wire2063, wire2062, wire2061, wire2060, wire2059, wire2058, wire2057, wire2056, wire2055, wire2054, wire2053, wire2052, wire2051, wire2050, wire2049, wire2048, wire2047, wire2046, wire2045, wire2044, wire2043, wire2042, wire2041, wire2040, wire2039, wire2038, wire2037, wire2036, wire2035, wire2034, wire2033, wire2032, wire2031, wire2030, wire2029, wire2028, wire2027, wire2026, wire2025, wire2024, wire2023, wire2022, wire2021, wire2020, wire2019, wire2018, wire2017, wire2016, wire2015, wire2014, wire2013, wire2012, wire2011, wire2010, wire2009, wire2008, wire2007, wire2006, wire2005, wire2004, wire2003, wire2002, wire2001, wire2000, wire1999, wire1998, wire1997, wire1996, wire1995, wire1994, wire1993, wire1992, wire1991, wire1990, wire1989, wire1988, wire1987, wire1986, wire1985, wire1984, wire1983, wire1982, wire1981, wire1980, wire1979, wire1978, wire1977, wire1976, wire1975, wire1974, wire1973, wire1972, wire1971, wire1970, wire1969, wire1968, wire1967, wire1966, wire1965, wire1964, wire1963, wire1962, wire1961, wire1960, wire1959, wire1958, wire1957, wire1956, wire1955, wire1954, wire1953, wire1952, wire1951, wire1950, wire1949, wire1948, wire1947, wire1946, wire1945, wire1944, wire1943, wire1942, wire1941, wire1940, wire1939, wire1938, wire1937, wire1936, wire1935, wire1934, wire1933, wire1932, wire1931, wire1930, wire1929, wire1928, wire1927, wire1926, wire1925, wire1924, wire1923, wire1922, wire1921, wire1920, wire1919, wire1918, wire1917, wire1916, wire1915, wire1914, wire1913, wire1912, wire1911, wire1910, wire1909, wire1908, wire1907, wire1906, wire1905, wire1904, wire1903, wire1902, wire1901, wire1900, wire1899, wire1898, wire1897, wire1896, wire1895, wire1894, wire1893, wire1892, wire1891, wire1890, wire1889, wire1888, wire1887, wire1886, wire1885, wire1884, wire1883, wire1882, wire1881, wire1880, wire1879, wire1878, wire1877, wire1876, wire1875, wire1874, wire1873, wire1872, wire1871, wire1870, wire1869, wire1868, wire1867, wire1866, wire1865, wire1864, wire1863, wire1862, wire1861, wire1860, wire1859, wire1858, wire1857, wire1856, wire1855, wire1854, wire1853, wire1852, wire1851, wire1850, wire1849, wire1848, wire1847, wire1846, wire1845, wire1844, wire1843, wire1842, wire1841, wire1840, wire1839, wire1838, wire1837, wire1836, wire1835, wire1834, wire1833, wire1832, wire1831, wire1830, wire1829, wire1828, wire1827, wire1826, wire1825, wire1824, wire1823, wire1822, wire1821, wire1820, wire1819, wire1818, wire1817, wire1816, wire1815, wire1814, wire1813, wire1812, wire1811, wire1810, wire1809, wire1808, wire1807, wire1806, wire1805, wire1804, wire1803, wire1802, wire1801, wire1800, wire1799, wire1798, wire1797, wire1796, wire1795, wire1794, wire1793, wire1792, wire1791, wire1790, wire1789, wire1788, wire1787, wire1786, wire1785, wire1784, wire1783, wire1782, wire1781, wire1780, wire1779, wire1778, wire1777, wire1776, wire1775, wire1774, wire1773, wire1772, wire1771, wire1770, wire1769, wire1768, wire1767, wire1766, wire1765, wire1764, wire1763, wire1762, wire1761, wire1760, wire1759, wire1758, wire1757, wire1756, wire1755, wire1754, wire1753, wire1752, wire1751, wire1750, wire1749, wire1748, wire1747, wire1746, wire1745, wire1744, wire1743, wire1742, wire1741, wire1740, wire1739, wire1738, wire1737, wire1736, wire1735, wire1734, wire1733, wire1732, wire1731, wire1730, wire1729, wire1728, wire1727, wire1726, wire1725, wire1724, wire1723, wire1722, wire1721, wire1720, wire1719, wire1718, wire1717, wire1716, wire1715, wire1714, wire1713, wire1712, wire1711, wire1710, wire1709, wire1708, wire1707, wire1706, wire1705, wire1704, wire1703, wire1702, wire1701, wire1700, wire1699, wire1698, wire1697, wire1696, wire1695, wire1694, wire1693, wire1692, wire1691, wire1690, wire1689, wire1688, wire1687, wire1686, wire1685, wire1684, wire1683, wire1682, wire1681, wire1680, wire1679, wire1678, wire1677, wire1676, wire1675, wire1674, wire1673, wire1672, wire1671, wire1670, wire1669, wire1668, wire1667, wire1666, wire1665, wire1664, wire1663, wire1662, wire1661, wire1660, wire1659, wire1658, wire1657, wire1656, wire1655, wire1654, wire1653, wire1652, wire1651, wire1650, wire1649, wire1648, wire1647, wire1646, wire1645, wire1644, wire1643, wire1642, wire1641, wire1640, wire1639, wire1638, wire1637, wire1636, wire1635, wire1634, wire1633, wire1632, wire1631, wire1630, wire1629, wire1628, wire1627, wire1626, wire1625, wire1624, wire1623, wire1622, wire1621, wire1620, wire1619, wire1618, wire1617, wire1616, wire1615, wire1614, wire1613, wire1612, wire1611, wire1610, wire1609, wire1608, wire1607, wire1606, wire1605, wire1604, wire1603, wire1602, wire1601, wire1600, wire1599, wire1598, wire1597, wire1596, wire1595, wire1594, wire1593, wire1592, wire1591, wire1590, wire1589, wire1588, wire1587, wire1586, wire1585, wire1584, wire1583, wire1582, wire1581, wire1580, wire1579, wire1578, wire1577, wire1576, wire1575, wire1574, wire1573, wire1572, wire1571, wire1570, wire1569, wire1568, wire1567, wire1566, wire1565, wire1564, wire1563, wire1562, wire1561, wire1560, wire1559, wire1558, wire1557, wire1556, wire1555, wire1554, wire1553, wire1552, wire1551, wire1550, wire1549, wire1548, wire1547, wire1546, wire1545, wire1544, wire1543, wire1542, wire1541, wire1540, wire1539, wire1538, wire1537, wire1536, wire1535, wire1534, wire1533, wire1532, wire1531, wire1530, wire1529, wire1528, wire1527, wire1526, wire1525, wire1524, wire1523, wire1522, wire1521, wire1520, wire1519, wire1518, wire1517, wire1516, wire1515, wire1514, wire1513, wire1512, wire1511, wire1510, wire1509, wire1508, wire1507, wire1506, wire1505, wire1504, wire1503, wire1502, wire1501, wire1500, wire1499, wire1498, wire1497, wire1496, wire1495, wire1494, wire1493, wire1492, wire1491, wire1490, wire1489, wire1488, wire1487, wire1486, wire1485, wire1484, wire1483, wire1482, wire1481, wire1480, wire1479, wire1478, wire1477, wire1476, wire1475, wire1474, wire1473, wire1472, wire1471, wire1470, wire1469, wire1468, wire1467, wire1466, wire1465, wire1464, wire1463, wire1462, wire1461, wire1460, wire1459, wire1458, wire1457, wire1456, wire1455, wire1454, wire1453, wire1452, wire1451, wire1450, wire1449, wire1448, wire1447, wire1446, wire1445, wire1444, wire1443, wire1442, wire1441, wire1440, wire1439, wire1438, wire1437, wire1436, wire1435, wire1434, wire1433, wire1432, wire1431, wire1430, wire1429, wire1428, wire1427, wire1426, wire1425, wire1424, wire1423, wire1422, wire1421, wire1420, wire1419, wire1418, wire1417, wire1416, wire1415, wire1414, wire1413, wire1412, wire1411, wire1410, wire1409, wire1408, wire1407, wire1406, wire1405, wire1404, wire1403, wire1402, wire1401, wire1400, wire1399, wire1398, wire1397, wire1396, wire1395, wire1394, wire1393, wire1392, wire1391, wire1390, wire1389, wire1388, wire1387, wire1386, wire1385, wire1384, wire1383, wire1382, wire1381, wire1380, wire1379, wire1378, wire1377, wire1376, wire1375, wire1374, wire1373, wire1372, wire1371, wire1370, wire1369, wire1368, wire1367, wire1366, wire1365, wire1364, wire1363, wire1362, wire1361, wire1360, wire1359, wire1358, wire1357, wire1356, wire1355, wire1354, wire1353, wire1352, wire1351, wire1350, wire1349, wire1348, wire1347, wire1346, wire1345, wire1344, wire1343, wire1342, wire1341, wire1340, wire1339, wire1338, wire1337, wire1336, wire1335, wire1334, wire1333, wire1332, wire1331, wire1330, wire1329, wire1328, wire1327, wire1326, wire1325, wire1324, wire1323, wire1322, wire1321, wire1320, wire1319, wire1318, wire1317, wire1316, wire1315, wire1314, wire1313, wire1312, wire1311, wire1310, wire1309, wire1308, wire1307, wire1306, wire1305, wire1304, wire1303, wire1302, wire1301, wire1300, wire1299, wire1298, wire1297, wire1296, wire1295, wire1294, wire1293, wire1292, wire1291, wire1290, wire1289, wire1288, wire1287, wire1286, wire1285, wire1284, wire1283, wire1282, wire1281, wire1280, wire1279, wire1278, wire1277, wire1276, wire1275, wire1274, wire1273, wire1272, wire1271, wire1270, wire1269, wire1268, wire1267, wire1266, wire1265, wire1264, wire1263, wire1262, wire1261, wire1260, wire1259, wire1258, wire1257, wire1256, wire1255, wire1254, wire1253, wire1252, wire1251, wire1250, wire1249, wire1248, wire1247, wire1246, wire1245, wire1244, wire1243, wire1242, wire1241, wire1240, wire1239, wire1238, wire1237, wire1236, wire1235, wire1234, wire1233, wire1232, wire1231, wire1230, wire1229, wire1228, wire1227, wire1226, wire1225, wire1224, wire1223, wire1222, wire1221, wire1220, wire1219, wire1218, wire1217, wire1216, wire1215, wire1214, wire1213, wire1212, wire1211, wire1210, wire1209, wire1208, wire1207, wire1206, wire1205, wire1204, wire1203, wire1202, wire1201, wire1200, wire1199, wire1198, wire1197, wire1196, wire1195, wire1194, wire1193, wire1192, wire1191, wire1190, wire1189, wire1188, wire1187, wire1186, wire1185, wire1184, wire1183, wire1182, wire1181, wire1180, wire1179, wire1178, wire1177, wire1176, wire1175, wire1174, wire1173, wire1172, wire1171, wire1170, wire1169, wire1168, wire1167, wire1166, wire1165, wire1164, wire1163, wire1162, wire1161, wire1160, wire1159, wire1158, wire1157, wire1156, wire1155, wire1154, wire1153, wire1152, wire1151, wire1150, wire1149, wire1148, wire1147, wire1146, wire1145, wire1144, wire1143, wire1142, wire1141, wire1140, wire1139, wire1138, wire1137, wire1136, wire1135, wire1134, wire1133, wire1132, wire1131, wire1130, wire1129, wire1128, wire1127, wire1126, wire1125, wire1124, wire1123, wire1122, wire1121, wire1120, wire1119, wire1118, wire1117, wire1116, wire1115, wire1114, wire1113, wire1112, wire1111, wire1110, wire1109, wire1108, wire1107, wire1106, wire1105, wire1104, wire1103, wire1102, wire1101, wire1100, wire1099, wire1098, wire1097, wire1096, wire1095, wire1094, wire1093, wire1092, wire1091, wire1090, wire1089, wire1088, wire1087, wire1086, wire1085, wire1084, wire1083, wire1082, wire1081, wire1080, wire1079, wire1078, wire1077, wire1076, wire1075, wire1074, wire1073, wire1072, wire1071, wire1070, wire1069, wire1068, wire1067, wire1066, wire1065, wire1064, wire1063, wire1062, wire1061, wire1060, wire1059, wire1058, wire1057, wire1056, wire1055, wire1054, wire1053, wire1052, wire1051, wire1050, wire1049, wire1048, wire1047, wire1046, wire1045, wire1044, wire1043, wire1042, wire1041, wire1040, wire1039, wire1038, wire1037, wire1036, wire1035, wire1034, wire1033, wire1032, wire1031, wire1030, wire1029, wire1028, wire1027, wire1026, wire1025, wire1024, wire1023, wire1022, wire1021, wire1020, wire1019, wire1018, wire1017, wire1016, wire1015, wire1014, wire1013, wire1012, wire1011, wire1010, wire1009, wire1008, wire1007, wire1006, wire1005, wire1004, wire1003, wire1002, wire1001, wire1000, wire999, wire998, wire997, wire996, wire995, wire994, wire993, wire992, wire991, wire990, wire989, wire988, wire987, wire986, wire985, wire984, wire983, wire982, wire981, wire980, wire979, wire978, wire977, wire976, wire975, wire974, wire973, wire972, wire971, wire970, wire969, wire968, wire967, wire966, wire965, wire964, wire963, wire962, wire961, wire960, wire959, wire958, wire957, wire956, wire955, wire954, wire953, wire952, wire951, wire950, wire949, wire948, wire947, wire946, wire945, wire944, wire943, wire942, wire941, wire940, wire939, wire938, wire937, wire936, wire935, wire934, wire933, wire932, wire931, wire930, wire929, wire928, wire927, wire926, wire925, wire924, wire923, wire922, wire921, wire920, wire919, wire918, wire917, wire916, wire915, wire914, wire913, wire912, wire911, wire910, wire909, wire908, wire907, wire906, wire905, wire904, wire903, wire902, wire901, wire900, wire899, wire898, wire897, wire896, wire895, wire894, wire893, wire892, wire891, wire890, wire889, wire888, wire887, wire886, wire885, wire884, wire883, wire882, wire881, wire880, wire879, wire878, wire877, wire876, wire875, wire874, wire873, wire872, wire871, wire870, wire869, wire868, wire867, wire866, wire865, wire864, wire863, wire862, wire861, wire860, wire859, wire858, wire857, wire856, wire855, wire854, wire853, wire852, wire851, wire850, wire849, wire848, wire847, wire846, wire845, wire844, wire843, wire842, wire841, wire840, wire839, wire838, wire837, wire836, wire835, wire834, wire833, wire832, wire831, wire830, wire829, wire828, wire827, wire826, wire825, wire824, wire823, wire822, wire821, wire820, wire819, wire818, wire817, wire816, wire815, wire814, wire813, wire812, wire811, wire810, wire809, wire808, wire807, wire806, wire805, wire804, wire803, wire802, wire801, wire800, wire799, wire798, wire797, wire796, wire795, wire794, wire793, wire792, wire791, wire790, wire789, wire788, wire787, wire786, wire785, wire784, wire783, wire782, wire781, wire780, wire779, wire778, wire777, wire776, wire775, wire774, wire773, wire772, wire771, wire770, wire769, wire768, wire767, wire766, wire765, wire764, wire763, wire762, wire761, wire760, wire759, wire758, wire757, wire756, wire755, wire754, wire753, wire752, wire751, wire750, wire749, wire748, wire747, wire746, wire745, wire744, wire743, wire742, wire741, wire740, wire739, wire738, wire737, wire736, wire735, wire734, wire733, wire732, wire731, wire730, wire729, wire728, wire727, wire726, wire725, wire724, wire723, wire722, wire721, wire720, wire719, wire718, wire717, wire716, wire715, wire714, wire713, wire712, wire711, wire710, wire709, wire708, wire707, wire706, wire705, wire704, wire703, wire702, wire701, wire700, wire699, wire698, wire697, wire696, wire695, wire694, wire693, wire692, wire691, wire690, wire689, wire688, wire687, wire686, wire685, wire684, wire683, wire682, wire681, wire680, wire679, wire678, wire677, wire676, wire675, wire674, wire673, wire672, wire671, wire670, wire669, wire668, wire667, wire666, wire665, wire664, wire663, wire662, wire661, wire660, wire659, wire658, wire657, wire656, wire655, wire654, wire653, wire652, wire651, wire650, wire649, wire648, wire647, wire646, wire645, wire644, wire643, wire642, wire641, wire640, wire639, wire638, wire637, wire636, wire635, wire634, wire633, wire632, wire631, wire630, wire629, wire628, wire627, wire626, wire625, wire624, wire623, wire622, wire621, wire620, wire619, wire618, wire617, wire616, wire615, wire614, wire613, wire612, wire611, wire610, wire609, wire608, wire607, wire606, wire605, wire604, wire603, wire602, wire601, wire600, wire599, wire598, wire597, wire596, wire595, wire594, wire593, wire592, wire591, wire590, wire589, wire588, wire587, wire586, wire585, wire584, wire583, wire582, wire581, wire580, wire579, wire578, wire577, wire576, wire575, wire574, wire573, wire572, wire571, wire570, wire569, wire568, wire567, wire566, wire565, wire564, wire563, wire562, wire561, wire560, wire559, wire558, wire557, wire556, wire555, wire554, wire553, wire552, wire551, wire550, wire549, wire548, wire547, wire546, wire545, wire544, wire543, wire542, wire541, wire540, wire539, wire538, wire537, wire536, wire535, wire534, wire533, wire532, wire531, wire530, wire529, wire528, wire527, wire526, wire525, wire524, wire523, wire522, wire521, wire520, wire519, wire518, wire517, wire516, wire515, wire514, wire513, wire512, wire511, wire510, wire509, wire508, wire507, wire506, wire505, wire504, wire503, wire502, wire501, wire500, wire499, wire498, wire497, wire496, wire495, wire494, wire493, wire492, wire491, wire490, wire489, wire488, wire487, wire486, wire485, wire484, wire483, wire482, wire481, wire480, wire479, wire478, wire477, wire476, wire475, wire474, wire473, wire472, wire471, wire470, wire469, wire468, wire467, wire466, wire465, wire464, wire463, wire462, wire461, wire460, wire459, wire458, wire457, wire456, wire455, wire454, wire453, wire452, wire451, wire450, wire449, wire448, wire447, wire446, wire445, wire444, wire443, wire442, wire441, wire440, wire439, wire438, wire437, wire436, wire435, wire434, wire433, wire432, wire431, wire430, wire429, wire428, wire427, wire426, wire425, wire424, wire423, wire422, wire421, wire420, wire419, wire418, wire417, wire416, wire415, wire414, wire413, wire412, wire411, wire410, wire409, wire408, wire407, wire406, wire405, wire404, wire403, wire402, wire401, wire400, wire399, wire398, wire397, wire396, wire395, wire394, wire393, wire392, wire391, wire390, wire389, wire388, wire387, wire386, wire385, wire384, wire383, wire382, wire381, wire380, wire379, wire378, wire377, wire376, wire375, wire374, wire373, wire372, wire371, wire370, wire369, wire368, wire367, wire366, wire365, wire364, wire363, wire362, wire361, wire360, wire359, wire358, wire357, wire356, wire355, wire354, wire353, wire352, wire351, wire350, wire349, wire348, wire347, wire346, wire345, wire344, wire343, wire342, wire341, wire340, wire339, wire338, wire337, wire336, wire335, wire334, wire333, wire332, wire331, wire330, wire329, wire328, wire327, wire326, wire325, wire324, wire323, wire322, wire321, wire320, wire319, wire318, wire317, wire316, wire315, wire314, wire313, wire312, wire311, wire310, wire309, wire308, wire307, wire306, wire305, wire304, wire303, wire302, wire301, wire300, wire299, wire298, wire297, wire296, wire295, wire294, wire293, wire292, wire291, wire290, wire289, wire288, wire287, wire286, wire285, wire284, wire283, wire282, wire281, wire280, wire279, wire278, wire277, wire276, wire275, wire274, wire273, wire272, wire271, wire270, wire269, wire268, wire267, wire266, wire265, wire264, wire263, wire262, wire261, wire260, wire259, wire258, wire257, wire256, wire255, wire254, wire253, wire252, wire251, wire250, wire249, wire248, wire247, wire246, wire245, wire244, wire243, wire242, wire241, wire240, wire239, wire238, wire237, wire236, wire235, wire234, wire233, wire232, wire231, wire230, wire229, wire228, wire227, wire226, wire225, wire224, wire223, wire222, wire221, wire220, wire219, wire218, wire217, wire216, wire215, wire214, wire213, wire212, wire211, wire210, wire209, wire208, wire207, wire206, wire205, wire204, wire203, wire202, wire201, wire200, wire199, wire198, wire197, wire196, wire195, wire194, wire193, wire192, wire191, wire190, wire189, wire188, wire187, wire186, wire185, wire184, wire183, wire182, wire181, wire180, wire179, wire178, wire177, wire176, wire175, wire174, wire173, wire172, wire171, wire170, wire169, wire168, wire167, wire166, wire165, wire164, wire163, wire162, wire161, wire160, wire159, wire158, wire157, wire156, wire155, wire154, wire153, wire152, wire151, wire150, wire149, wire148, wire147, wire146, wire145, wire144, wire143, wire142, wire141, wire140, wire139, wire138, wire137, wire136, wire135, wire134, wire133, wire132, wire131, wire130, wire129, wire128, wire127, wire126, wire125, wire124, wire123, wire122, wire121, wire120, wire119, wire118, wire117, wire116, wire115, wire114, wire113, wire112, wire111, wire110, wire109, wire108, wire107, wire106, wire105, wire104, wire103, wire102, wire101, wire100, wire99, wire98, wire97, wire96, wire95, wire94, wire93, wire92, wire91, wire90, wire89, wire88, wire87, wire86, wire85, wire84, wire83, wire82, wire81, wire80, wire79, wire78, wire77, wire76, wire75, wire74, wire73, wire72, wire71, wire70, wire69, wire68, wire67, wire66, wire65, wire64, wire63, wire62, wire61, wire60, wire59, wire58, wire57, wire56, wire55, wire54, wire53, wire52, wire51, wire50, wire49, wire48, wire47, wire46, wire45, wire44, wire43, wire42, wire41, wire40, wire39, wire38, wire37, wire36, wire35, wire34, wire33, wire32, wire31, wire30, wire29, wire28, wire27, wire26, wire25, wire24, wire23, wire22, wire21, wire20, wire19, wire18, wire17, wire16, wire15, wire14, wire13, wire12, wire11, wire10, wire9, wire8, wire7, wire6, wire5, wire4, wire3, wire2, wire1, wire0};

    muxnm_tristate #(4096, 8) mxt1(.in(data_concat), .sel(weq_concat) ,.out(out));
endmodule
