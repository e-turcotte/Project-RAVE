module select_length(
    input wire [11:0] sel,
    output wire [7:0] out
);
    wire [3071:0] data;
    length_data ld(.out(data));
    wire [383:0] sel_out;
    select_signal s0(.sel(sel), .out(sel_out));
    muxnm_tristate #(384, 8) mxt1(.in(data), .sel(sel_out) ,.out(out));

endmodule

module select_signal(
    input wire [11:0] sel,
    output wire [383:0] out
);
    wire [11:0] buffered_input;
    bufferH1024_nb$ #(12) buff(.in(sel), .out(buffered_input));
    equaln #(12) e0(.a(buffered_input), .b(12'b000000000001), .eq(weq0));
    equaln #(12) e1(.a(buffered_input), .b(12'b010000000001), .eq(weq1));
    equaln #(12) e2(.a(buffered_input), .b(12'b100000000001), .eq(weq2));
    equaln #(12) e3(.a(buffered_input), .b(12'b110000000001), .eq(weq3));
    equaln #(12) e4(.a(buffered_input), .b(12'b001000000001), .eq(weq4));
    equaln #(12) e5(.a(buffered_input), .b(12'b011000000001), .eq(weq5));
    equaln #(12) e6(.a(buffered_input), .b(12'b101000000001), .eq(weq6));
    equaln #(12) e7(.a(buffered_input), .b(12'b111000000001), .eq(weq7));
    equaln #(12) e8(.a(buffered_input), .b(12'b000100000001), .eq(weq8));
    equaln #(12) e9(.a(buffered_input), .b(12'b010100000001), .eq(weq9));
    equaln #(12) e10(.a(buffered_input), .b(12'b100100000001), .eq(weq10));
    equaln #(12) e11(.a(buffered_input), .b(12'b110100000001), .eq(weq11));
    equaln #(12) e12(.a(buffered_input), .b(12'b001100000001), .eq(weq12));
    equaln #(12) e13(.a(buffered_input), .b(12'b011100000001), .eq(weq13));
    equaln #(12) e14(.a(buffered_input), .b(12'b101100000001), .eq(weq14));
    equaln #(12) e15(.a(buffered_input), .b(12'b111100000001), .eq(weq15));
    equaln #(12) e16(.a(buffered_input), .b(12'b000001000001), .eq(weq16));
    equaln #(12) e17(.a(buffered_input), .b(12'b010001000001), .eq(weq17));
    equaln #(12) e18(.a(buffered_input), .b(12'b100001000001), .eq(weq18));
    equaln #(12) e19(.a(buffered_input), .b(12'b110001000001), .eq(weq19));
    equaln #(12) e20(.a(buffered_input), .b(12'b001001000001), .eq(weq20));
    equaln #(12) e21(.a(buffered_input), .b(12'b011001000001), .eq(weq21));
    equaln #(12) e22(.a(buffered_input), .b(12'b101001000001), .eq(weq22));
    equaln #(12) e23(.a(buffered_input), .b(12'b111001000001), .eq(weq23));
    equaln #(12) e24(.a(buffered_input), .b(12'b000101000001), .eq(weq24));
    equaln #(12) e25(.a(buffered_input), .b(12'b010101000001), .eq(weq25));
    equaln #(12) e26(.a(buffered_input), .b(12'b100101000001), .eq(weq26));
    equaln #(12) e27(.a(buffered_input), .b(12'b110101000001), .eq(weq27));
    equaln #(12) e28(.a(buffered_input), .b(12'b001101000001), .eq(weq28));
    equaln #(12) e29(.a(buffered_input), .b(12'b011101000001), .eq(weq29));
    equaln #(12) e30(.a(buffered_input), .b(12'b101101000001), .eq(weq30));
    equaln #(12) e31(.a(buffered_input), .b(12'b111101000001), .eq(weq31));
    equaln #(12) e32(.a(buffered_input), .b(12'b000010000001), .eq(weq32));
    equaln #(12) e33(.a(buffered_input), .b(12'b010010000001), .eq(weq33));
    equaln #(12) e34(.a(buffered_input), .b(12'b100010000001), .eq(weq34));
    equaln #(12) e35(.a(buffered_input), .b(12'b110010000001), .eq(weq35));
    equaln #(12) e36(.a(buffered_input), .b(12'b001010000001), .eq(weq36));
    equaln #(12) e37(.a(buffered_input), .b(12'b011010000001), .eq(weq37));
    equaln #(12) e38(.a(buffered_input), .b(12'b101010000001), .eq(weq38));
    equaln #(12) e39(.a(buffered_input), .b(12'b111010000001), .eq(weq39));
    equaln #(12) e40(.a(buffered_input), .b(12'b000110000001), .eq(weq40));
    equaln #(12) e41(.a(buffered_input), .b(12'b010110000001), .eq(weq41));
    equaln #(12) e42(.a(buffered_input), .b(12'b100110000001), .eq(weq42));
    equaln #(12) e43(.a(buffered_input), .b(12'b110110000001), .eq(weq43));
    equaln #(12) e44(.a(buffered_input), .b(12'b001110000001), .eq(weq44));
    equaln #(12) e45(.a(buffered_input), .b(12'b011110000001), .eq(weq45));
    equaln #(12) e46(.a(buffered_input), .b(12'b101110000001), .eq(weq46));
    equaln #(12) e47(.a(buffered_input), .b(12'b111110000001), .eq(weq47));
    equaln #(12) e48(.a(buffered_input), .b(12'b000011000001), .eq(weq48));
    equaln #(12) e49(.a(buffered_input), .b(12'b010011000001), .eq(weq49));
    equaln #(12) e50(.a(buffered_input), .b(12'b100011000001), .eq(weq50));
    equaln #(12) e51(.a(buffered_input), .b(12'b110011000001), .eq(weq51));
    equaln #(12) e52(.a(buffered_input), .b(12'b001011000001), .eq(weq52));
    equaln #(12) e53(.a(buffered_input), .b(12'b011011000001), .eq(weq53));
    equaln #(12) e54(.a(buffered_input), .b(12'b101011000001), .eq(weq54));
    equaln #(12) e55(.a(buffered_input), .b(12'b111011000001), .eq(weq55));
    equaln #(12) e56(.a(buffered_input), .b(12'b000111000001), .eq(weq56));
    equaln #(12) e57(.a(buffered_input), .b(12'b010111000001), .eq(weq57));
    equaln #(12) e58(.a(buffered_input), .b(12'b100111000001), .eq(weq58));
    equaln #(12) e59(.a(buffered_input), .b(12'b110111000001), .eq(weq59));
    equaln #(12) e60(.a(buffered_input), .b(12'b001111000001), .eq(weq60));
    equaln #(12) e61(.a(buffered_input), .b(12'b011111000001), .eq(weq61));
    equaln #(12) e62(.a(buffered_input), .b(12'b101111000001), .eq(weq62));
    equaln #(12) e63(.a(buffered_input), .b(12'b111111000001), .eq(weq63));
    equaln #(12) e64(.a(buffered_input), .b(12'b000000000010), .eq(weq64));
    equaln #(12) e65(.a(buffered_input), .b(12'b010000000010), .eq(weq65));
    equaln #(12) e66(.a(buffered_input), .b(12'b100000000010), .eq(weq66));
    equaln #(12) e67(.a(buffered_input), .b(12'b110000000010), .eq(weq67));
    equaln #(12) e68(.a(buffered_input), .b(12'b001000000010), .eq(weq68));
    equaln #(12) e69(.a(buffered_input), .b(12'b011000000010), .eq(weq69));
    equaln #(12) e70(.a(buffered_input), .b(12'b101000000010), .eq(weq70));
    equaln #(12) e71(.a(buffered_input), .b(12'b111000000010), .eq(weq71));
    equaln #(12) e72(.a(buffered_input), .b(12'b000100000010), .eq(weq72));
    equaln #(12) e73(.a(buffered_input), .b(12'b010100000010), .eq(weq73));
    equaln #(12) e74(.a(buffered_input), .b(12'b100100000010), .eq(weq74));
    equaln #(12) e75(.a(buffered_input), .b(12'b110100000010), .eq(weq75));
    equaln #(12) e76(.a(buffered_input), .b(12'b001100000010), .eq(weq76));
    equaln #(12) e77(.a(buffered_input), .b(12'b011100000010), .eq(weq77));
    equaln #(12) e78(.a(buffered_input), .b(12'b101100000010), .eq(weq78));
    equaln #(12) e79(.a(buffered_input), .b(12'b111100000010), .eq(weq79));
    equaln #(12) e80(.a(buffered_input), .b(12'b000001000010), .eq(weq80));
    equaln #(12) e81(.a(buffered_input), .b(12'b010001000010), .eq(weq81));
    equaln #(12) e82(.a(buffered_input), .b(12'b100001000010), .eq(weq82));
    equaln #(12) e83(.a(buffered_input), .b(12'b110001000010), .eq(weq83));
    equaln #(12) e84(.a(buffered_input), .b(12'b001001000010), .eq(weq84));
    equaln #(12) e85(.a(buffered_input), .b(12'b011001000010), .eq(weq85));
    equaln #(12) e86(.a(buffered_input), .b(12'b101001000010), .eq(weq86));
    equaln #(12) e87(.a(buffered_input), .b(12'b111001000010), .eq(weq87));
    equaln #(12) e88(.a(buffered_input), .b(12'b000101000010), .eq(weq88));
    equaln #(12) e89(.a(buffered_input), .b(12'b010101000010), .eq(weq89));
    equaln #(12) e90(.a(buffered_input), .b(12'b100101000010), .eq(weq90));
    equaln #(12) e91(.a(buffered_input), .b(12'b110101000010), .eq(weq91));
    equaln #(12) e92(.a(buffered_input), .b(12'b001101000010), .eq(weq92));
    equaln #(12) e93(.a(buffered_input), .b(12'b011101000010), .eq(weq93));
    equaln #(12) e94(.a(buffered_input), .b(12'b101101000010), .eq(weq94));
    equaln #(12) e95(.a(buffered_input), .b(12'b111101000010), .eq(weq95));
    equaln #(12) e96(.a(buffered_input), .b(12'b000010000010), .eq(weq96));
    equaln #(12) e97(.a(buffered_input), .b(12'b010010000010), .eq(weq97));
    equaln #(12) e98(.a(buffered_input), .b(12'b100010000010), .eq(weq98));
    equaln #(12) e99(.a(buffered_input), .b(12'b110010000010), .eq(weq99));
    equaln #(12) e100(.a(buffered_input), .b(12'b001010000010), .eq(weq100));
    equaln #(12) e101(.a(buffered_input), .b(12'b011010000010), .eq(weq101));
    equaln #(12) e102(.a(buffered_input), .b(12'b101010000010), .eq(weq102));
    equaln #(12) e103(.a(buffered_input), .b(12'b111010000010), .eq(weq103));
    equaln #(12) e104(.a(buffered_input), .b(12'b000110000010), .eq(weq104));
    equaln #(12) e105(.a(buffered_input), .b(12'b010110000010), .eq(weq105));
    equaln #(12) e106(.a(buffered_input), .b(12'b100110000010), .eq(weq106));
    equaln #(12) e107(.a(buffered_input), .b(12'b110110000010), .eq(weq107));
    equaln #(12) e108(.a(buffered_input), .b(12'b001110000010), .eq(weq108));
    equaln #(12) e109(.a(buffered_input), .b(12'b011110000010), .eq(weq109));
    equaln #(12) e110(.a(buffered_input), .b(12'b101110000010), .eq(weq110));
    equaln #(12) e111(.a(buffered_input), .b(12'b111110000010), .eq(weq111));
    equaln #(12) e112(.a(buffered_input), .b(12'b000011000010), .eq(weq112));
    equaln #(12) e113(.a(buffered_input), .b(12'b010011000010), .eq(weq113));
    equaln #(12) e114(.a(buffered_input), .b(12'b100011000010), .eq(weq114));
    equaln #(12) e115(.a(buffered_input), .b(12'b110011000010), .eq(weq115));
    equaln #(12) e116(.a(buffered_input), .b(12'b001011000010), .eq(weq116));
    equaln #(12) e117(.a(buffered_input), .b(12'b011011000010), .eq(weq117));
    equaln #(12) e118(.a(buffered_input), .b(12'b101011000010), .eq(weq118));
    equaln #(12) e119(.a(buffered_input), .b(12'b111011000010), .eq(weq119));
    equaln #(12) e120(.a(buffered_input), .b(12'b000111000010), .eq(weq120));
    equaln #(12) e121(.a(buffered_input), .b(12'b010111000010), .eq(weq121));
    equaln #(12) e122(.a(buffered_input), .b(12'b100111000010), .eq(weq122));
    equaln #(12) e123(.a(buffered_input), .b(12'b110111000010), .eq(weq123));
    equaln #(12) e124(.a(buffered_input), .b(12'b001111000010), .eq(weq124));
    equaln #(12) e125(.a(buffered_input), .b(12'b011111000010), .eq(weq125));
    equaln #(12) e126(.a(buffered_input), .b(12'b101111000010), .eq(weq126));
    equaln #(12) e127(.a(buffered_input), .b(12'b111111000010), .eq(weq127));
    equaln #(12) e128(.a(buffered_input), .b(12'b000000000100), .eq(weq128));
    equaln #(12) e129(.a(buffered_input), .b(12'b010000000100), .eq(weq129));
    equaln #(12) e130(.a(buffered_input), .b(12'b100000000100), .eq(weq130));
    equaln #(12) e131(.a(buffered_input), .b(12'b110000000100), .eq(weq131));
    equaln #(12) e132(.a(buffered_input), .b(12'b001000000100), .eq(weq132));
    equaln #(12) e133(.a(buffered_input), .b(12'b011000000100), .eq(weq133));
    equaln #(12) e134(.a(buffered_input), .b(12'b101000000100), .eq(weq134));
    equaln #(12) e135(.a(buffered_input), .b(12'b111000000100), .eq(weq135));
    equaln #(12) e136(.a(buffered_input), .b(12'b000100000100), .eq(weq136));
    equaln #(12) e137(.a(buffered_input), .b(12'b010100000100), .eq(weq137));
    equaln #(12) e138(.a(buffered_input), .b(12'b100100000100), .eq(weq138));
    equaln #(12) e139(.a(buffered_input), .b(12'b110100000100), .eq(weq139));
    equaln #(12) e140(.a(buffered_input), .b(12'b001100000100), .eq(weq140));
    equaln #(12) e141(.a(buffered_input), .b(12'b011100000100), .eq(weq141));
    equaln #(12) e142(.a(buffered_input), .b(12'b101100000100), .eq(weq142));
    equaln #(12) e143(.a(buffered_input), .b(12'b111100000100), .eq(weq143));
    equaln #(12) e144(.a(buffered_input), .b(12'b000001000100), .eq(weq144));
    equaln #(12) e145(.a(buffered_input), .b(12'b010001000100), .eq(weq145));
    equaln #(12) e146(.a(buffered_input), .b(12'b100001000100), .eq(weq146));
    equaln #(12) e147(.a(buffered_input), .b(12'b110001000100), .eq(weq147));
    equaln #(12) e148(.a(buffered_input), .b(12'b001001000100), .eq(weq148));
    equaln #(12) e149(.a(buffered_input), .b(12'b011001000100), .eq(weq149));
    equaln #(12) e150(.a(buffered_input), .b(12'b101001000100), .eq(weq150));
    equaln #(12) e151(.a(buffered_input), .b(12'b111001000100), .eq(weq151));
    equaln #(12) e152(.a(buffered_input), .b(12'b000101000100), .eq(weq152));
    equaln #(12) e153(.a(buffered_input), .b(12'b010101000100), .eq(weq153));
    equaln #(12) e154(.a(buffered_input), .b(12'b100101000100), .eq(weq154));
    equaln #(12) e155(.a(buffered_input), .b(12'b110101000100), .eq(weq155));
    equaln #(12) e156(.a(buffered_input), .b(12'b001101000100), .eq(weq156));
    equaln #(12) e157(.a(buffered_input), .b(12'b011101000100), .eq(weq157));
    equaln #(12) e158(.a(buffered_input), .b(12'b101101000100), .eq(weq158));
    equaln #(12) e159(.a(buffered_input), .b(12'b111101000100), .eq(weq159));
    equaln #(12) e160(.a(buffered_input), .b(12'b000010000100), .eq(weq160));
    equaln #(12) e161(.a(buffered_input), .b(12'b010010000100), .eq(weq161));
    equaln #(12) e162(.a(buffered_input), .b(12'b100010000100), .eq(weq162));
    equaln #(12) e163(.a(buffered_input), .b(12'b110010000100), .eq(weq163));
    equaln #(12) e164(.a(buffered_input), .b(12'b001010000100), .eq(weq164));
    equaln #(12) e165(.a(buffered_input), .b(12'b011010000100), .eq(weq165));
    equaln #(12) e166(.a(buffered_input), .b(12'b101010000100), .eq(weq166));
    equaln #(12) e167(.a(buffered_input), .b(12'b111010000100), .eq(weq167));
    equaln #(12) e168(.a(buffered_input), .b(12'b000110000100), .eq(weq168));
    equaln #(12) e169(.a(buffered_input), .b(12'b010110000100), .eq(weq169));
    equaln #(12) e170(.a(buffered_input), .b(12'b100110000100), .eq(weq170));
    equaln #(12) e171(.a(buffered_input), .b(12'b110110000100), .eq(weq171));
    equaln #(12) e172(.a(buffered_input), .b(12'b001110000100), .eq(weq172));
    equaln #(12) e173(.a(buffered_input), .b(12'b011110000100), .eq(weq173));
    equaln #(12) e174(.a(buffered_input), .b(12'b101110000100), .eq(weq174));
    equaln #(12) e175(.a(buffered_input), .b(12'b111110000100), .eq(weq175));
    equaln #(12) e176(.a(buffered_input), .b(12'b000011000100), .eq(weq176));
    equaln #(12) e177(.a(buffered_input), .b(12'b010011000100), .eq(weq177));
    equaln #(12) e178(.a(buffered_input), .b(12'b100011000100), .eq(weq178));
    equaln #(12) e179(.a(buffered_input), .b(12'b110011000100), .eq(weq179));
    equaln #(12) e180(.a(buffered_input), .b(12'b001011000100), .eq(weq180));
    equaln #(12) e181(.a(buffered_input), .b(12'b011011000100), .eq(weq181));
    equaln #(12) e182(.a(buffered_input), .b(12'b101011000100), .eq(weq182));
    equaln #(12) e183(.a(buffered_input), .b(12'b111011000100), .eq(weq183));
    equaln #(12) e184(.a(buffered_input), .b(12'b000111000100), .eq(weq184));
    equaln #(12) e185(.a(buffered_input), .b(12'b010111000100), .eq(weq185));
    equaln #(12) e186(.a(buffered_input), .b(12'b100111000100), .eq(weq186));
    equaln #(12) e187(.a(buffered_input), .b(12'b110111000100), .eq(weq187));
    equaln #(12) e188(.a(buffered_input), .b(12'b001111000100), .eq(weq188));
    equaln #(12) e189(.a(buffered_input), .b(12'b011111000100), .eq(weq189));
    equaln #(12) e190(.a(buffered_input), .b(12'b101111000100), .eq(weq190));
    equaln #(12) e191(.a(buffered_input), .b(12'b111111000100), .eq(weq191));
    equaln #(12) e192(.a(buffered_input), .b(12'b000000001000), .eq(weq192));
    equaln #(12) e193(.a(buffered_input), .b(12'b010000001000), .eq(weq193));
    equaln #(12) e194(.a(buffered_input), .b(12'b100000001000), .eq(weq194));
    equaln #(12) e195(.a(buffered_input), .b(12'b110000001000), .eq(weq195));
    equaln #(12) e196(.a(buffered_input), .b(12'b001000001000), .eq(weq196));
    equaln #(12) e197(.a(buffered_input), .b(12'b011000001000), .eq(weq197));
    equaln #(12) e198(.a(buffered_input), .b(12'b101000001000), .eq(weq198));
    equaln #(12) e199(.a(buffered_input), .b(12'b111000001000), .eq(weq199));
    equaln #(12) e200(.a(buffered_input), .b(12'b000100001000), .eq(weq200));
    equaln #(12) e201(.a(buffered_input), .b(12'b010100001000), .eq(weq201));
    equaln #(12) e202(.a(buffered_input), .b(12'b100100001000), .eq(weq202));
    equaln #(12) e203(.a(buffered_input), .b(12'b110100001000), .eq(weq203));
    equaln #(12) e204(.a(buffered_input), .b(12'b001100001000), .eq(weq204));
    equaln #(12) e205(.a(buffered_input), .b(12'b011100001000), .eq(weq205));
    equaln #(12) e206(.a(buffered_input), .b(12'b101100001000), .eq(weq206));
    equaln #(12) e207(.a(buffered_input), .b(12'b111100001000), .eq(weq207));
    equaln #(12) e208(.a(buffered_input), .b(12'b000001001000), .eq(weq208));
    equaln #(12) e209(.a(buffered_input), .b(12'b010001001000), .eq(weq209));
    equaln #(12) e210(.a(buffered_input), .b(12'b100001001000), .eq(weq210));
    equaln #(12) e211(.a(buffered_input), .b(12'b110001001000), .eq(weq211));
    equaln #(12) e212(.a(buffered_input), .b(12'b001001001000), .eq(weq212));
    equaln #(12) e213(.a(buffered_input), .b(12'b011001001000), .eq(weq213));
    equaln #(12) e214(.a(buffered_input), .b(12'b101001001000), .eq(weq214));
    equaln #(12) e215(.a(buffered_input), .b(12'b111001001000), .eq(weq215));
    equaln #(12) e216(.a(buffered_input), .b(12'b000101001000), .eq(weq216));
    equaln #(12) e217(.a(buffered_input), .b(12'b010101001000), .eq(weq217));
    equaln #(12) e218(.a(buffered_input), .b(12'b100101001000), .eq(weq218));
    equaln #(12) e219(.a(buffered_input), .b(12'b110101001000), .eq(weq219));
    equaln #(12) e220(.a(buffered_input), .b(12'b001101001000), .eq(weq220));
    equaln #(12) e221(.a(buffered_input), .b(12'b011101001000), .eq(weq221));
    equaln #(12) e222(.a(buffered_input), .b(12'b101101001000), .eq(weq222));
    equaln #(12) e223(.a(buffered_input), .b(12'b111101001000), .eq(weq223));
    equaln #(12) e224(.a(buffered_input), .b(12'b000010001000), .eq(weq224));
    equaln #(12) e225(.a(buffered_input), .b(12'b010010001000), .eq(weq225));
    equaln #(12) e226(.a(buffered_input), .b(12'b100010001000), .eq(weq226));
    equaln #(12) e227(.a(buffered_input), .b(12'b110010001000), .eq(weq227));
    equaln #(12) e228(.a(buffered_input), .b(12'b001010001000), .eq(weq228));
    equaln #(12) e229(.a(buffered_input), .b(12'b011010001000), .eq(weq229));
    equaln #(12) e230(.a(buffered_input), .b(12'b101010001000), .eq(weq230));
    equaln #(12) e231(.a(buffered_input), .b(12'b111010001000), .eq(weq231));
    equaln #(12) e232(.a(buffered_input), .b(12'b000110001000), .eq(weq232));
    equaln #(12) e233(.a(buffered_input), .b(12'b010110001000), .eq(weq233));
    equaln #(12) e234(.a(buffered_input), .b(12'b100110001000), .eq(weq234));
    equaln #(12) e235(.a(buffered_input), .b(12'b110110001000), .eq(weq235));
    equaln #(12) e236(.a(buffered_input), .b(12'b001110001000), .eq(weq236));
    equaln #(12) e237(.a(buffered_input), .b(12'b011110001000), .eq(weq237));
    equaln #(12) e238(.a(buffered_input), .b(12'b101110001000), .eq(weq238));
    equaln #(12) e239(.a(buffered_input), .b(12'b111110001000), .eq(weq239));
    equaln #(12) e240(.a(buffered_input), .b(12'b000011001000), .eq(weq240));
    equaln #(12) e241(.a(buffered_input), .b(12'b010011001000), .eq(weq241));
    equaln #(12) e242(.a(buffered_input), .b(12'b100011001000), .eq(weq242));
    equaln #(12) e243(.a(buffered_input), .b(12'b110011001000), .eq(weq243));
    equaln #(12) e244(.a(buffered_input), .b(12'b001011001000), .eq(weq244));
    equaln #(12) e245(.a(buffered_input), .b(12'b011011001000), .eq(weq245));
    equaln #(12) e246(.a(buffered_input), .b(12'b101011001000), .eq(weq246));
    equaln #(12) e247(.a(buffered_input), .b(12'b111011001000), .eq(weq247));
    equaln #(12) e248(.a(buffered_input), .b(12'b000111001000), .eq(weq248));
    equaln #(12) e249(.a(buffered_input), .b(12'b010111001000), .eq(weq249));
    equaln #(12) e250(.a(buffered_input), .b(12'b100111001000), .eq(weq250));
    equaln #(12) e251(.a(buffered_input), .b(12'b110111001000), .eq(weq251));
    equaln #(12) e252(.a(buffered_input), .b(12'b001111001000), .eq(weq252));
    equaln #(12) e253(.a(buffered_input), .b(12'b011111001000), .eq(weq253));
    equaln #(12) e254(.a(buffered_input), .b(12'b101111001000), .eq(weq254));
    equaln #(12) e255(.a(buffered_input), .b(12'b111111001000), .eq(weq255));
    equaln #(12) e256(.a(buffered_input), .b(12'b000000010000), .eq(weq256));
    equaln #(12) e257(.a(buffered_input), .b(12'b010000010000), .eq(weq257));
    equaln #(12) e258(.a(buffered_input), .b(12'b100000010000), .eq(weq258));
    equaln #(12) e259(.a(buffered_input), .b(12'b110000010000), .eq(weq259));
    equaln #(12) e260(.a(buffered_input), .b(12'b001000010000), .eq(weq260));
    equaln #(12) e261(.a(buffered_input), .b(12'b011000010000), .eq(weq261));
    equaln #(12) e262(.a(buffered_input), .b(12'b101000010000), .eq(weq262));
    equaln #(12) e263(.a(buffered_input), .b(12'b111000010000), .eq(weq263));
    equaln #(12) e264(.a(buffered_input), .b(12'b000100010000), .eq(weq264));
    equaln #(12) e265(.a(buffered_input), .b(12'b010100010000), .eq(weq265));
    equaln #(12) e266(.a(buffered_input), .b(12'b100100010000), .eq(weq266));
    equaln #(12) e267(.a(buffered_input), .b(12'b110100010000), .eq(weq267));
    equaln #(12) e268(.a(buffered_input), .b(12'b001100010000), .eq(weq268));
    equaln #(12) e269(.a(buffered_input), .b(12'b011100010000), .eq(weq269));
    equaln #(12) e270(.a(buffered_input), .b(12'b101100010000), .eq(weq270));
    equaln #(12) e271(.a(buffered_input), .b(12'b111100010000), .eq(weq271));
    equaln #(12) e272(.a(buffered_input), .b(12'b000001010000), .eq(weq272));
    equaln #(12) e273(.a(buffered_input), .b(12'b010001010000), .eq(weq273));
    equaln #(12) e274(.a(buffered_input), .b(12'b100001010000), .eq(weq274));
    equaln #(12) e275(.a(buffered_input), .b(12'b110001010000), .eq(weq275));
    equaln #(12) e276(.a(buffered_input), .b(12'b001001010000), .eq(weq276));
    equaln #(12) e277(.a(buffered_input), .b(12'b011001010000), .eq(weq277));
    equaln #(12) e278(.a(buffered_input), .b(12'b101001010000), .eq(weq278));
    equaln #(12) e279(.a(buffered_input), .b(12'b111001010000), .eq(weq279));
    equaln #(12) e280(.a(buffered_input), .b(12'b000101010000), .eq(weq280));
    equaln #(12) e281(.a(buffered_input), .b(12'b010101010000), .eq(weq281));
    equaln #(12) e282(.a(buffered_input), .b(12'b100101010000), .eq(weq282));
    equaln #(12) e283(.a(buffered_input), .b(12'b110101010000), .eq(weq283));
    equaln #(12) e284(.a(buffered_input), .b(12'b001101010000), .eq(weq284));
    equaln #(12) e285(.a(buffered_input), .b(12'b011101010000), .eq(weq285));
    equaln #(12) e286(.a(buffered_input), .b(12'b101101010000), .eq(weq286));
    equaln #(12) e287(.a(buffered_input), .b(12'b111101010000), .eq(weq287));
    equaln #(12) e288(.a(buffered_input), .b(12'b000010010000), .eq(weq288));
    equaln #(12) e289(.a(buffered_input), .b(12'b010010010000), .eq(weq289));
    equaln #(12) e290(.a(buffered_input), .b(12'b100010010000), .eq(weq290));
    equaln #(12) e291(.a(buffered_input), .b(12'b110010010000), .eq(weq291));
    equaln #(12) e292(.a(buffered_input), .b(12'b001010010000), .eq(weq292));
    equaln #(12) e293(.a(buffered_input), .b(12'b011010010000), .eq(weq293));
    equaln #(12) e294(.a(buffered_input), .b(12'b101010010000), .eq(weq294));
    equaln #(12) e295(.a(buffered_input), .b(12'b111010010000), .eq(weq295));
    equaln #(12) e296(.a(buffered_input), .b(12'b000110010000), .eq(weq296));
    equaln #(12) e297(.a(buffered_input), .b(12'b010110010000), .eq(weq297));
    equaln #(12) e298(.a(buffered_input), .b(12'b100110010000), .eq(weq298));
    equaln #(12) e299(.a(buffered_input), .b(12'b110110010000), .eq(weq299));
    equaln #(12) e300(.a(buffered_input), .b(12'b001110010000), .eq(weq300));
    equaln #(12) e301(.a(buffered_input), .b(12'b011110010000), .eq(weq301));
    equaln #(12) e302(.a(buffered_input), .b(12'b101110010000), .eq(weq302));
    equaln #(12) e303(.a(buffered_input), .b(12'b111110010000), .eq(weq303));
    equaln #(12) e304(.a(buffered_input), .b(12'b000011010000), .eq(weq304));
    equaln #(12) e305(.a(buffered_input), .b(12'b010011010000), .eq(weq305));
    equaln #(12) e306(.a(buffered_input), .b(12'b100011010000), .eq(weq306));
    equaln #(12) e307(.a(buffered_input), .b(12'b110011010000), .eq(weq307));
    equaln #(12) e308(.a(buffered_input), .b(12'b001011010000), .eq(weq308));
    equaln #(12) e309(.a(buffered_input), .b(12'b011011010000), .eq(weq309));
    equaln #(12) e310(.a(buffered_input), .b(12'b101011010000), .eq(weq310));
    equaln #(12) e311(.a(buffered_input), .b(12'b111011010000), .eq(weq311));
    equaln #(12) e312(.a(buffered_input), .b(12'b000111010000), .eq(weq312));
    equaln #(12) e313(.a(buffered_input), .b(12'b010111010000), .eq(weq313));
    equaln #(12) e314(.a(buffered_input), .b(12'b100111010000), .eq(weq314));
    equaln #(12) e315(.a(buffered_input), .b(12'b110111010000), .eq(weq315));
    equaln #(12) e316(.a(buffered_input), .b(12'b001111010000), .eq(weq316));
    equaln #(12) e317(.a(buffered_input), .b(12'b011111010000), .eq(weq317));
    equaln #(12) e318(.a(buffered_input), .b(12'b101111010000), .eq(weq318));
    equaln #(12) e319(.a(buffered_input), .b(12'b111111010000), .eq(weq319));
    equaln #(12) e320(.a(buffered_input), .b(12'b000000100000), .eq(weq320));
    equaln #(12) e321(.a(buffered_input), .b(12'b010000100000), .eq(weq321));
    equaln #(12) e322(.a(buffered_input), .b(12'b100000100000), .eq(weq322));
    equaln #(12) e323(.a(buffered_input), .b(12'b110000100000), .eq(weq323));
    equaln #(12) e324(.a(buffered_input), .b(12'b001000100000), .eq(weq324));
    equaln #(12) e325(.a(buffered_input), .b(12'b011000100000), .eq(weq325));
    equaln #(12) e326(.a(buffered_input), .b(12'b101000100000), .eq(weq326));
    equaln #(12) e327(.a(buffered_input), .b(12'b111000100000), .eq(weq327));
    equaln #(12) e328(.a(buffered_input), .b(12'b000100100000), .eq(weq328));
    equaln #(12) e329(.a(buffered_input), .b(12'b010100100000), .eq(weq329));
    equaln #(12) e330(.a(buffered_input), .b(12'b100100100000), .eq(weq330));
    equaln #(12) e331(.a(buffered_input), .b(12'b110100100000), .eq(weq331));
    equaln #(12) e332(.a(buffered_input), .b(12'b001100100000), .eq(weq332));
    equaln #(12) e333(.a(buffered_input), .b(12'b011100100000), .eq(weq333));
    equaln #(12) e334(.a(buffered_input), .b(12'b101100100000), .eq(weq334));
    equaln #(12) e335(.a(buffered_input), .b(12'b111100100000), .eq(weq335));
    equaln #(12) e336(.a(buffered_input), .b(12'b000001100000), .eq(weq336));
    equaln #(12) e337(.a(buffered_input), .b(12'b010001100000), .eq(weq337));
    equaln #(12) e338(.a(buffered_input), .b(12'b100001100000), .eq(weq338));
    equaln #(12) e339(.a(buffered_input), .b(12'b110001100000), .eq(weq339));
    equaln #(12) e340(.a(buffered_input), .b(12'b001001100000), .eq(weq340));
    equaln #(12) e341(.a(buffered_input), .b(12'b011001100000), .eq(weq341));
    equaln #(12) e342(.a(buffered_input), .b(12'b101001100000), .eq(weq342));
    equaln #(12) e343(.a(buffered_input), .b(12'b111001100000), .eq(weq343));
    equaln #(12) e344(.a(buffered_input), .b(12'b000101100000), .eq(weq344));
    equaln #(12) e345(.a(buffered_input), .b(12'b010101100000), .eq(weq345));
    equaln #(12) e346(.a(buffered_input), .b(12'b100101100000), .eq(weq346));
    equaln #(12) e347(.a(buffered_input), .b(12'b110101100000), .eq(weq347));
    equaln #(12) e348(.a(buffered_input), .b(12'b001101100000), .eq(weq348));
    equaln #(12) e349(.a(buffered_input), .b(12'b011101100000), .eq(weq349));
    equaln #(12) e350(.a(buffered_input), .b(12'b101101100000), .eq(weq350));
    equaln #(12) e351(.a(buffered_input), .b(12'b111101100000), .eq(weq351));
    equaln #(12) e352(.a(buffered_input), .b(12'b000010100000), .eq(weq352));
    equaln #(12) e353(.a(buffered_input), .b(12'b010010100000), .eq(weq353));
    equaln #(12) e354(.a(buffered_input), .b(12'b100010100000), .eq(weq354));
    equaln #(12) e355(.a(buffered_input), .b(12'b110010100000), .eq(weq355));
    equaln #(12) e356(.a(buffered_input), .b(12'b001010100000), .eq(weq356));
    equaln #(12) e357(.a(buffered_input), .b(12'b011010100000), .eq(weq357));
    equaln #(12) e358(.a(buffered_input), .b(12'b101010100000), .eq(weq358));
    equaln #(12) e359(.a(buffered_input), .b(12'b111010100000), .eq(weq359));
    equaln #(12) e360(.a(buffered_input), .b(12'b000110100000), .eq(weq360));
    equaln #(12) e361(.a(buffered_input), .b(12'b010110100000), .eq(weq361));
    equaln #(12) e362(.a(buffered_input), .b(12'b100110100000), .eq(weq362));
    equaln #(12) e363(.a(buffered_input), .b(12'b110110100000), .eq(weq363));
    equaln #(12) e364(.a(buffered_input), .b(12'b001110100000), .eq(weq364));
    equaln #(12) e365(.a(buffered_input), .b(12'b011110100000), .eq(weq365));
    equaln #(12) e366(.a(buffered_input), .b(12'b101110100000), .eq(weq366));
    equaln #(12) e367(.a(buffered_input), .b(12'b111110100000), .eq(weq367));
    equaln #(12) e368(.a(buffered_input), .b(12'b000011100000), .eq(weq368));
    equaln #(12) e369(.a(buffered_input), .b(12'b010011100000), .eq(weq369));
    equaln #(12) e370(.a(buffered_input), .b(12'b100011100000), .eq(weq370));
    equaln #(12) e371(.a(buffered_input), .b(12'b110011100000), .eq(weq371));
    equaln #(12) e372(.a(buffered_input), .b(12'b001011100000), .eq(weq372));
    equaln #(12) e373(.a(buffered_input), .b(12'b011011100000), .eq(weq373));
    equaln #(12) e374(.a(buffered_input), .b(12'b101011100000), .eq(weq374));
    equaln #(12) e375(.a(buffered_input), .b(12'b111011100000), .eq(weq375));
    equaln #(12) e376(.a(buffered_input), .b(12'b000111100000), .eq(weq376));
    equaln #(12) e377(.a(buffered_input), .b(12'b010111100000), .eq(weq377));
    equaln #(12) e378(.a(buffered_input), .b(12'b100111100000), .eq(weq378));
    equaln #(12) e379(.a(buffered_input), .b(12'b110111100000), .eq(weq379));
    equaln #(12) e380(.a(buffered_input), .b(12'b001111100000), .eq(weq380));
    equaln #(12) e381(.a(buffered_input), .b(12'b011111100000), .eq(weq381));
    equaln #(12) e382(.a(buffered_input), .b(12'b101111100000), .eq(weq382));
    equaln #(12) e383(.a(buffered_input), .b(12'b111111100000), .eq(weq383));
    assign out = {weq383, weq382, weq381, weq380, weq379, weq378, weq377, weq376, weq375, weq374, weq373, weq372, weq371, weq370, weq369, weq368, weq367, weq366, weq365, weq364, weq363, weq362, weq361, weq360, weq359, weq358, weq357, weq356, weq355, weq354, weq353, weq352, weq351, weq350, weq349, weq348, weq347, weq346, weq345, weq344, weq343, weq342, weq341, weq340, weq339, weq338, weq337, weq336, weq335, weq334, weq333, weq332, weq331, weq330, weq329, weq328, weq327, weq326, weq325, weq324, weq323, weq322, weq321, weq320, weq319, weq318, weq317, weq316, weq315, weq314, weq313, weq312, weq311, weq310, weq309, weq308, weq307, weq306, weq305, weq304, weq303, weq302, weq301, weq300, weq299, weq298, weq297, weq296, weq295, weq294, weq293, weq292, weq291, weq290, weq289, weq288, weq287, weq286, weq285, weq284, weq283, weq282, weq281, weq280, weq279, weq278, weq277, weq276, weq275, weq274, weq273, weq272, weq271, weq270, weq269, weq268, weq267, weq266, weq265, weq264, weq263, weq262, weq261, weq260, weq259, weq258, weq257, weq256, weq255, weq254, weq253, weq252, weq251, weq250, weq249, weq248, weq247, weq246, weq245, weq244, weq243, weq242, weq241, weq240, weq239, weq238, weq237, weq236, weq235, weq234, weq233, weq232, weq231, weq230, weq229, weq228, weq227, weq226, weq225, weq224, weq223, weq222, weq221, weq220, weq219, weq218, weq217, weq216, weq215, weq214, weq213, weq212, weq211, weq210, weq209, weq208, weq207, weq206, weq205, weq204, weq203, weq202, weq201, weq200, weq199, weq198, weq197, weq196, weq195, weq194, weq193, weq192, weq191, weq190, weq189, weq188, weq187, weq186, weq185, weq184, weq183, weq182, weq181, weq180, weq179, weq178, weq177, weq176, weq175, weq174, weq173, weq172, weq171, weq170, weq169, weq168, weq167, weq166, weq165, weq164, weq163, weq162, weq161, weq160, weq159, weq158, weq157, weq156, weq155, weq154, weq153, weq152, weq151, weq150, weq149, weq148, weq147, weq146, weq145, weq144, weq143, weq142, weq141, weq140, weq139, weq138, weq137, weq136, weq135, weq134, weq133, weq132, weq131, weq130, weq129, weq128, weq127, weq126, weq125, weq124, weq123, weq122, weq121, weq120, weq119, weq118, weq117, weq116, weq115, weq114, weq113, weq112, weq111, weq110, weq109, weq108, weq107, weq106, weq105, weq104, weq103, weq102, weq101, weq100, weq99, weq98, weq97, weq96, weq95, weq94, weq93, weq92, weq91, weq90, weq89, weq88, weq87, weq86, weq85, weq84, weq83, weq82, weq81, weq80, weq79, weq78, weq77, weq76, weq75, weq74, weq73, weq72, weq71, weq70, weq69, weq68, weq67, weq66, weq65, weq64, weq63, weq62, weq61, weq60, weq59, weq58, weq57, weq56, weq55, weq54, weq53, weq52, weq51, weq50, weq49, weq48, weq47, weq46, weq45, weq44, weq43, weq42, weq41, weq40, weq39, weq38, weq37, weq36, weq35, weq34, weq33, weq32, weq31, weq30, weq29, weq28, weq27, weq26, weq25, weq24, weq23, weq22, weq21, weq20, weq19, weq18, weq17, weq16, weq15, weq14, weq13, weq12, weq11, weq10, weq9, weq8, weq7, weq6, weq5, weq4, weq3, weq2, weq1, weq0};


endmodule