module eflags_t();

endmodule