module TOP;

    reg [3:0] recvB, grantB, ackB;
    reg bus_clk, clr;
    wire [72:0] BUS;
    wire [3:0] freeB, relB, reqB;

    pmem_TOP pm(.recvB(recvB), .grantB(grantB), .ackB(ackB), .bus_clk(bus_clk), .clr(clr),
                .BUS(BUS), .freeB(freeB), .relB(relB), .reqB(reqB));

    initial begin
        $readmemh("initfiles/pmem_b0c0d0.init", pm.banks[0].bnk.bank_slices[0].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c0d1.init", pm.banks[0].bnk.bank_slices[0].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c0d2.init", pm.banks[0].bnk.bank_slices[0].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c0d3.init", pm.banks[0].bnk.bank_slices[0].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c1d0.init", pm.banks[0].bnk.bank_slices[1].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c1d1.init", pm.banks[0].bnk.bank_slices[1].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c1d2.init", pm.banks[0].bnk.bank_slices[1].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c1d3.init", pm.banks[0].bnk.bank_slices[1].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c2d0.init", pm.banks[0].bnk.bank_slices[2].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c2d1.init", pm.banks[0].bnk.bank_slices[2].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c2d2.init", pm.banks[0].bnk.bank_slices[2].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c2d3.init", pm.banks[0].bnk.bank_slices[2].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c3d0.init", pm.banks[0].bnk.bank_slices[3].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c3d1.init", pm.banks[0].bnk.bank_slices[3].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c3d2.init", pm.banks[0].bnk.bank_slices[3].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c3d3.init", pm.banks[0].bnk.bank_slices[3].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c4d0.init", pm.banks[0].bnk.bank_slices[4].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c4d1.init", pm.banks[0].bnk.bank_slices[4].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c4d2.init", pm.banks[0].bnk.bank_slices[4].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c4d3.init", pm.banks[0].bnk.bank_slices[4].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c5d0.init", pm.banks[0].bnk.bank_slices[5].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c5d1.init", pm.banks[0].bnk.bank_slices[5].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c5d2.init", pm.banks[0].bnk.bank_slices[5].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c5d3.init", pm.banks[0].bnk.bank_slices[5].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c6d0.init", pm.banks[0].bnk.bank_slices[6].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c6d1.init", pm.banks[0].bnk.bank_slices[6].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c6d2.init", pm.banks[0].bnk.bank_slices[6].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c6d3.init", pm.banks[0].bnk.bank_slices[6].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c7d0.init", pm.banks[0].bnk.bank_slices[7].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c7d1.init", pm.banks[0].bnk.bank_slices[7].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c7d2.init", pm.banks[0].bnk.bank_slices[7].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c7d3.init", pm.banks[0].bnk.bank_slices[7].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c8d0.init", pm.banks[0].bnk.bank_slices[8].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c8d1.init", pm.banks[0].bnk.bank_slices[8].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c8d2.init", pm.banks[0].bnk.bank_slices[8].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c8d3.init", pm.banks[0].bnk.bank_slices[8].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c9d0.init", pm.banks[0].bnk.bank_slices[9].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c9d1.init", pm.banks[0].bnk.bank_slices[9].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c9d2.init", pm.banks[0].bnk.bank_slices[9].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c9d3.init", pm.banks[0].bnk.bank_slices[9].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c10d0.init", pm.banks[0].bnk.bank_slices[10].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c10d1.init", pm.banks[0].bnk.bank_slices[10].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c10d2.init", pm.banks[0].bnk.bank_slices[10].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c10d3.init", pm.banks[0].bnk.bank_slices[10].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c11d0.init", pm.banks[0].bnk.bank_slices[11].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c11d1.init", pm.banks[0].bnk.bank_slices[11].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c11d2.init", pm.banks[0].bnk.bank_slices[11].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c11d3.init", pm.banks[0].bnk.bank_slices[11].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c12d0.init", pm.banks[0].bnk.bank_slices[12].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c12d1.init", pm.banks[0].bnk.bank_slices[12].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c12d2.init", pm.banks[0].bnk.bank_slices[12].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c12d3.init", pm.banks[0].bnk.bank_slices[12].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c13d0.init", pm.banks[0].bnk.bank_slices[13].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c13d1.init", pm.banks[0].bnk.bank_slices[13].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c13d2.init", pm.banks[0].bnk.bank_slices[13].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c13d3.init", pm.banks[0].bnk.bank_slices[13].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c14d0.init", pm.banks[0].bnk.bank_slices[14].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c14d1.init", pm.banks[0].bnk.bank_slices[14].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c14d2.init", pm.banks[0].bnk.bank_slices[14].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c14d3.init", pm.banks[0].bnk.bank_slices[14].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b0c15d0.init", pm.banks[0].bnk.bank_slices[15].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b0c15d1.init", pm.banks[0].bnk.bank_slices[15].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b0c15d2.init", pm.banks[0].bnk.bank_slices[15].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b0c15d3.init", pm.banks[0].bnk.bank_slices[15].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c0d0.init", pm.banks[1].bnk.bank_slices[0].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c0d1.init", pm.banks[1].bnk.bank_slices[0].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c0d2.init", pm.banks[1].bnk.bank_slices[0].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c0d3.init", pm.banks[1].bnk.bank_slices[0].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c1d0.init", pm.banks[1].bnk.bank_slices[1].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c1d1.init", pm.banks[1].bnk.bank_slices[1].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c1d2.init", pm.banks[1].bnk.bank_slices[1].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c1d3.init", pm.banks[1].bnk.bank_slices[1].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c2d0.init", pm.banks[1].bnk.bank_slices[2].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c2d1.init", pm.banks[1].bnk.bank_slices[2].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c2d2.init", pm.banks[1].bnk.bank_slices[2].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c2d3.init", pm.banks[1].bnk.bank_slices[2].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c3d0.init", pm.banks[1].bnk.bank_slices[3].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c3d1.init", pm.banks[1].bnk.bank_slices[3].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c3d2.init", pm.banks[1].bnk.bank_slices[3].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c3d3.init", pm.banks[1].bnk.bank_slices[3].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c4d0.init", pm.banks[1].bnk.bank_slices[4].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c4d1.init", pm.banks[1].bnk.bank_slices[4].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c4d2.init", pm.banks[1].bnk.bank_slices[4].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c4d3.init", pm.banks[1].bnk.bank_slices[4].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c5d0.init", pm.banks[1].bnk.bank_slices[5].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c5d1.init", pm.banks[1].bnk.bank_slices[5].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c5d2.init", pm.banks[1].bnk.bank_slices[5].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c5d3.init", pm.banks[1].bnk.bank_slices[5].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c6d0.init", pm.banks[1].bnk.bank_slices[6].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c6d1.init", pm.banks[1].bnk.bank_slices[6].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c6d2.init", pm.banks[1].bnk.bank_slices[6].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c6d3.init", pm.banks[1].bnk.bank_slices[6].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c7d0.init", pm.banks[1].bnk.bank_slices[7].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c7d1.init", pm.banks[1].bnk.bank_slices[7].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c7d2.init", pm.banks[1].bnk.bank_slices[7].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c7d3.init", pm.banks[1].bnk.bank_slices[7].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c8d0.init", pm.banks[1].bnk.bank_slices[8].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c8d1.init", pm.banks[1].bnk.bank_slices[8].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c8d2.init", pm.banks[1].bnk.bank_slices[8].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c8d3.init", pm.banks[1].bnk.bank_slices[8].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c9d0.init", pm.banks[1].bnk.bank_slices[9].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c9d1.init", pm.banks[1].bnk.bank_slices[9].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c9d2.init", pm.banks[1].bnk.bank_slices[9].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c9d3.init", pm.banks[1].bnk.bank_slices[9].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c10d0.init", pm.banks[1].bnk.bank_slices[10].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c10d1.init", pm.banks[1].bnk.bank_slices[10].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c10d2.init", pm.banks[1].bnk.bank_slices[10].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c10d3.init", pm.banks[1].bnk.bank_slices[10].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c11d0.init", pm.banks[1].bnk.bank_slices[11].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c11d1.init", pm.banks[1].bnk.bank_slices[11].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c11d2.init", pm.banks[1].bnk.bank_slices[11].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c11d3.init", pm.banks[1].bnk.bank_slices[11].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c12d0.init", pm.banks[1].bnk.bank_slices[12].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c12d1.init", pm.banks[1].bnk.bank_slices[12].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c12d2.init", pm.banks[1].bnk.bank_slices[12].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c12d3.init", pm.banks[1].bnk.bank_slices[12].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c13d0.init", pm.banks[1].bnk.bank_slices[13].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c13d1.init", pm.banks[1].bnk.bank_slices[13].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c13d2.init", pm.banks[1].bnk.bank_slices[13].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c13d3.init", pm.banks[1].bnk.bank_slices[13].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c14d0.init", pm.banks[1].bnk.bank_slices[14].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c14d1.init", pm.banks[1].bnk.bank_slices[14].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c14d2.init", pm.banks[1].bnk.bank_slices[14].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c14d3.init", pm.banks[1].bnk.bank_slices[14].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b1c15d0.init", pm.banks[1].bnk.bank_slices[15].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b1c15d1.init", pm.banks[1].bnk.bank_slices[15].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b1c15d2.init", pm.banks[1].bnk.bank_slices[15].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b1c15d3.init", pm.banks[1].bnk.bank_slices[15].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c0d0.init", pm.banks[2].bnk.bank_slices[0].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c0d1.init", pm.banks[2].bnk.bank_slices[0].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c0d2.init", pm.banks[2].bnk.bank_slices[0].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c0d3.init", pm.banks[2].bnk.bank_slices[0].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c1d0.init", pm.banks[2].bnk.bank_slices[1].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c1d1.init", pm.banks[2].bnk.bank_slices[1].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c1d2.init", pm.banks[2].bnk.bank_slices[1].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c1d3.init", pm.banks[2].bnk.bank_slices[1].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c2d0.init", pm.banks[2].bnk.bank_slices[2].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c2d1.init", pm.banks[2].bnk.bank_slices[2].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c2d2.init", pm.banks[2].bnk.bank_slices[2].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c2d3.init", pm.banks[2].bnk.bank_slices[2].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c3d0.init", pm.banks[2].bnk.bank_slices[3].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c3d1.init", pm.banks[2].bnk.bank_slices[3].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c3d2.init", pm.banks[2].bnk.bank_slices[3].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c3d3.init", pm.banks[2].bnk.bank_slices[3].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c4d0.init", pm.banks[2].bnk.bank_slices[4].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c4d1.init", pm.banks[2].bnk.bank_slices[4].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c4d2.init", pm.banks[2].bnk.bank_slices[4].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c4d3.init", pm.banks[2].bnk.bank_slices[4].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c5d0.init", pm.banks[2].bnk.bank_slices[5].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c5d1.init", pm.banks[2].bnk.bank_slices[5].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c5d2.init", pm.banks[2].bnk.bank_slices[5].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c5d3.init", pm.banks[2].bnk.bank_slices[5].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c6d0.init", pm.banks[2].bnk.bank_slices[6].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c6d1.init", pm.banks[2].bnk.bank_slices[6].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c6d2.init", pm.banks[2].bnk.bank_slices[6].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c6d3.init", pm.banks[2].bnk.bank_slices[6].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c7d0.init", pm.banks[2].bnk.bank_slices[7].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c7d1.init", pm.banks[2].bnk.bank_slices[7].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c7d2.init", pm.banks[2].bnk.bank_slices[7].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c7d3.init", pm.banks[2].bnk.bank_slices[7].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c8d0.init", pm.banks[2].bnk.bank_slices[8].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c8d1.init", pm.banks[2].bnk.bank_slices[8].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c8d2.init", pm.banks[2].bnk.bank_slices[8].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c8d3.init", pm.banks[2].bnk.bank_slices[8].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c9d0.init", pm.banks[2].bnk.bank_slices[9].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c9d1.init", pm.banks[2].bnk.bank_slices[9].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c9d2.init", pm.banks[2].bnk.bank_slices[9].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c9d3.init", pm.banks[2].bnk.bank_slices[9].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c10d0.init", pm.banks[2].bnk.bank_slices[10].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c10d1.init", pm.banks[2].bnk.bank_slices[10].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c10d2.init", pm.banks[2].bnk.bank_slices[10].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c10d3.init", pm.banks[2].bnk.bank_slices[10].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c11d0.init", pm.banks[2].bnk.bank_slices[11].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c11d1.init", pm.banks[2].bnk.bank_slices[11].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c11d2.init", pm.banks[2].bnk.bank_slices[11].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c11d3.init", pm.banks[2].bnk.bank_slices[11].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c12d0.init", pm.banks[2].bnk.bank_slices[12].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c12d1.init", pm.banks[2].bnk.bank_slices[12].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c12d2.init", pm.banks[2].bnk.bank_slices[12].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c12d3.init", pm.banks[2].bnk.bank_slices[12].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c13d0.init", pm.banks[2].bnk.bank_slices[13].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c13d1.init", pm.banks[2].bnk.bank_slices[13].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c13d2.init", pm.banks[2].bnk.bank_slices[13].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c13d3.init", pm.banks[2].bnk.bank_slices[13].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c14d0.init", pm.banks[2].bnk.bank_slices[14].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c14d1.init", pm.banks[2].bnk.bank_slices[14].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c14d2.init", pm.banks[2].bnk.bank_slices[14].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c14d3.init", pm.banks[2].bnk.bank_slices[14].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b2c15d0.init", pm.banks[2].bnk.bank_slices[15].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b2c15d1.init", pm.banks[2].bnk.bank_slices[15].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b2c15d2.init", pm.banks[2].bnk.bank_slices[15].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b2c15d3.init", pm.banks[2].bnk.bank_slices[15].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c0d0.init", pm.banks[3].bnk.bank_slices[0].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c0d1.init", pm.banks[3].bnk.bank_slices[0].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c0d2.init", pm.banks[3].bnk.bank_slices[0].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c0d3.init", pm.banks[3].bnk.bank_slices[0].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c1d0.init", pm.banks[3].bnk.bank_slices[1].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c1d1.init", pm.banks[3].bnk.bank_slices[1].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c1d2.init", pm.banks[3].bnk.bank_slices[1].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c1d3.init", pm.banks[3].bnk.bank_slices[1].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c2d0.init", pm.banks[3].bnk.bank_slices[2].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c2d1.init", pm.banks[3].bnk.bank_slices[2].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c2d2.init", pm.banks[3].bnk.bank_slices[2].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c2d3.init", pm.banks[3].bnk.bank_slices[2].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c3d0.init", pm.banks[3].bnk.bank_slices[3].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c3d1.init", pm.banks[3].bnk.bank_slices[3].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c3d2.init", pm.banks[3].bnk.bank_slices[3].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c3d3.init", pm.banks[3].bnk.bank_slices[3].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c4d0.init", pm.banks[3].bnk.bank_slices[4].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c4d1.init", pm.banks[3].bnk.bank_slices[4].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c4d2.init", pm.banks[3].bnk.bank_slices[4].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c4d3.init", pm.banks[3].bnk.bank_slices[4].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c5d0.init", pm.banks[3].bnk.bank_slices[5].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c5d1.init", pm.banks[3].bnk.bank_slices[5].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c5d2.init", pm.banks[3].bnk.bank_slices[5].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c5d3.init", pm.banks[3].bnk.bank_slices[5].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c6d0.init", pm.banks[3].bnk.bank_slices[6].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c6d1.init", pm.banks[3].bnk.bank_slices[6].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c6d2.init", pm.banks[3].bnk.bank_slices[6].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c6d3.init", pm.banks[3].bnk.bank_slices[6].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c7d0.init", pm.banks[3].bnk.bank_slices[7].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c7d1.init", pm.banks[3].bnk.bank_slices[7].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c7d2.init", pm.banks[3].bnk.bank_slices[7].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c7d3.init", pm.banks[3].bnk.bank_slices[7].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c8d0.init", pm.banks[3].bnk.bank_slices[8].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c8d1.init", pm.banks[3].bnk.bank_slices[8].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c8d2.init", pm.banks[3].bnk.bank_slices[8].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c8d3.init", pm.banks[3].bnk.bank_slices[8].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c9d0.init", pm.banks[3].bnk.bank_slices[9].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c9d1.init", pm.banks[3].bnk.bank_slices[9].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c9d2.init", pm.banks[3].bnk.bank_slices[9].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c9d3.init", pm.banks[3].bnk.bank_slices[9].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c10d0.init", pm.banks[3].bnk.bank_slices[10].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c10d1.init", pm.banks[3].bnk.bank_slices[10].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c10d2.init", pm.banks[3].bnk.bank_slices[10].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c10d3.init", pm.banks[3].bnk.bank_slices[10].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c11d0.init", pm.banks[3].bnk.bank_slices[11].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c11d1.init", pm.banks[3].bnk.bank_slices[11].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c11d2.init", pm.banks[3].bnk.bank_slices[11].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c11d3.init", pm.banks[3].bnk.bank_slices[11].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c12d0.init", pm.banks[3].bnk.bank_slices[12].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c12d1.init", pm.banks[3].bnk.bank_slices[12].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c12d2.init", pm.banks[3].bnk.bank_slices[12].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c12d3.init", pm.banks[3].bnk.bank_slices[12].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c13d0.init", pm.banks[3].bnk.bank_slices[13].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c13d1.init", pm.banks[3].bnk.bank_slices[13].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c13d2.init", pm.banks[3].bnk.bank_slices[13].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c13d3.init", pm.banks[3].bnk.bank_slices[13].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c14d0.init", pm.banks[3].bnk.bank_slices[14].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c14d1.init", pm.banks[3].bnk.bank_slices[14].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c14d2.init", pm.banks[3].bnk.bank_slices[14].dram.cells[2].sram.mem);
        $readmemh("initfiles/pmem_b3c14d3.init", pm.banks[3].bnk.bank_slices[14].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c15d0.init", pm.banks[3].bnk.bank_slices[15].dram.cells[0].sram.mem);
        $readmemh("initfiles/pmem_b3c15d1.init", pm.banks[3].bnk.bank_slices[15].dram.cells[1].sram.mem);
        $readmemh("initfiles/pmem_b3c15d3.init", pm.banks[3].bnk.bank_slices[15].dram.cells[3].sram.mem);
        $readmemh("initfiles/pmem_b3c15d2.init", pm.banks[3].bnk.bank_slices[15].dram.cells[2].sram.mem);
    end

endmodule