module TOP();
    localparam CYCLE_TIME = 12.0;
    
    integer file;
    reg clk;
    integer cycle_number; //TODO
    
    initial begin
        file = $fopen("debug.out", "w");
        clk = 1'b1;
        cycle_number = 0;
        forever #(CYCLE_TIME / 2.0) clk = ~clk;
    end

    //TODO: TLB Initializations
    reg [19:0] VP_0, VP_1, VP_2, VP_3, VP_4, VP_5, VP_6, VP_7;
	reg [19:0] PF_0, PF_1, PF_2, PF_3, PF_4, PF_5, PF_6, PF_7;
	reg [7:0] entry_v;
	reg [7:0] entry_P;
	reg [7:0] entry_RW;
    reg [7:0] entry_PCD;
	reg [159:0] VP, PF; //concats of VP_7 to VP_0 and PF_7 to PF_0

    //TODO: Core initializations:
    reg global_reset;
    reg global_set;

    //Pipeline: FETCH1 -> FETCH2 -> DECODE -> RrAg -> MEM -> EX -> WB

    //  IMPORTANT NOTES:
    //   -  notation for latche wires: <signal.name>_<stage.prev>_<stage.next>_latch_<in/out>
    //      where <in> is the input to the latch (output of stage.prev) and <out> is the output 
    //      from the latch (input of stage.next)

    ///////////////////////////////////////////////////////////
    // Outputs from Rr/Ag that go into the RrAg_MEM_latch:  //  
    //////////////////////////////////////////////////////////
    
    wire         valid_RrAg_MEM_latch_in, stall_RrAg_MEM_latch_in;
    wire [1:0]   opsize_RrAg_MEM_latch_in;
    wire [31:0]  mem_addr1_RrAg_MEM_latch_in, mem_addr2_RrAg_MEM_latch_in, mem_addr1_end_RrAg_MEM_latch_in, mem_addr2_end_RrAg_MEM_latch_in;
    wire [63:0]  reg1_RrAg_MEM_latch_in, reg2_RrAg_MEM_latch_in, reg3_RrAg_MEM_latch_in, reg4_RrAg_MEM_latch_in;
    wire [127:0] ptc_r1_RrAg_MEM_latch_in, ptc_r2_RrAg_MEM_latch_in, ptc_r3_RrAg_MEM_latch_in, ptc_r4_RrAg_MEM_latch_in;
    wire [2:0]   reg1_orig_RrAg_MEM_latch_in, reg2_orig_RrAg_MEM_latch_in, reg3_orig_RrAg_MEM_latch_in, reg4_orig_RrAg_MEM_latch_in;
    wire [15:0]  seg1_RrAg_MEM_latch_in, seg2_RrAg_MEM_latch_in, seg3_RrAg_MEM_latch_in, seg4_RrAg_MEM_latch_in;
    wire [31:0]  ptc_s1_RrAg_MEM_latch_in, ptc_s2_RrAg_MEM_latch_in, ptc_s3_RrAg_MEM_latch_in, ptc_s4_RrAg_MEM_latch_in;
    wire [2:0]   seg1_orig_RrAg_MEM_latch_in, seg2_orig_RrAg_MEM_latch_in, seg3_orig_RrAg_MEM_latch_in, seg4_orig_RrAg_MEM_latch_in;
    wire [6:0]   inst_ptcid_RrAg_MEM_latch_in;
    wire [12:0]  op1_out_RrAg_MEM_latch_in, op2_out_RrAg_MEM_latch_in, op3_out_RrAg_MEM_latch_in, op4_out_RrAg_MEM_latch_in;
    wire [12:0]  dest1_out_RrAg_MEM_latch_in, dest2_out_RrAg_MEM_latch_in, dest3_out_RrAg_MEM_latch_in, dest4_out_RrAg_MEM_latch_in;
    wire         res1_ld_out_RrAg_MEM_latch_in, res2_ld_out_RrAg_MEM_latch_in, res3_ld_out_RrAg_MEM_latch_in, res4_ld_out_RrAg_MEM_latch_in;
    wire [31:0]  rep_num_RrAg_MEM_latch_in;
    wire [4:0]   aluk_out_RrAg_MEM_latch_in;
    wire [2:0]   mux_adder_out_RrAg_MEM_latch_in;
    wire         mux_and_int_out_RrAg_MEM_latch_in, mux_shift_out_RrAg_MEM_latch_in;
    wire [36:0]  p_op_out_RrAg_MEM_latch_in;
    wire [17:0]  fmask_out_RrAg_MEM_latch_in;
    wire [1:0]   conditionals_out_RrAg_MEM_latch_in;
    wire         is_br_out_RrAg_MEM_latch_in, is_fp_out_RrAg_MEM_latch_in;
    wire [47:0]  imm_out_RrAg_MEM_latch_in;
    wire [1:0]   mem1_rw_out_RrAg_MEM_latch_in, mem2_rw_out_RrAg_MEM_latch_in;
    wire [31:0]  eip_out_RrAg_MEM_latch_in;
    wire         IE_out_RrAg_MEM_latch_in;
    wire [3:0]   IE_type_out_RrAg_MEM_latch_in;
    wire [31:0]  BR_pred_target_out_RrAg_MEM_latch_in;
    wire         BR_pred_T_NT_out_RrAg_MEM_latch_in;
    
    ///////////////////////////////////////////////////////////
    //   Outputs from RrAg_MEM_latch that go into the MEM:  //  
    //////////////////////////////////////////////////////////

    wire         valid_RrAg_MEM_latch_out, stall_RrAg_MEM_latch_out;
    wire [1:0]   opsize_RrAg_MEM_latch_out;
    wire [31:0]  mem_addr1_RrAg_MEM_latch_out, mem_addr2_RrAg_MEM_latch_out, mem_addr1_end_RrAg_MEM_latch_out, mem_addr2_end_RrAg_MEM_latch_out;
    wire [63:0]  reg1_RrAg_MEM_latch_out, reg2_RrAg_MEM_latch_out, reg3_RrAg_MEM_latch_out, reg4_RrAg_MEM_latch_out;
    wire [127:0] ptc_r1_RrAg_MEM_latch_out, ptc_r2_RrAg_MEM_latch_out, ptc_r3_RrAg_MEM_latch_out, ptc_r4_RrAg_MEM_latch_out;
    wire [2:0]   reg1_orig_RrAg_MEM_latch_out, reg2_orig_RrAg_MEM_latch_out, reg3_orig_RrAg_MEM_latch_out, reg4_orig_RrAg_MEM_latch_out;
    wire [15:0]  seg1_RrAg_MEM_latch_out, seg2_RrAg_MEM_latch_out, seg3_RrAg_MEM_latch_out, seg4_RrAg_MEM_latch_out;
    wire [31:0]  ptc_s1_RrAg_MEM_latch_out, ptc_s2_RrAg_MEM_latch_out, ptc_s3_RrAg_MEM_latch_out, ptc_s4_RrAg_MEM_latch_out;
    wire [2:0]   seg1_orig_RrAg_MEM_latch_out, seg2_orig_RrAg_MEM_latch_out, seg3_orig_RrAg_MEM_latch_out, seg4_orig_RrAg_MEM_latch_out;
    wire [6:0]   inst_ptcid_RrAg_MEM_latch_out;
    wire [12:0]  op1_RrAg_MEM_latch_out, op2_RrAg_MEM_latch_out, op3_RrAg_MEM_latch_out, op4_RrAg_MEM_latch_out;
    wire [12:0]  dest1_RrAg_MEM_latch_out, dest2_RrAg_MEM_latch_out, dest3_RrAg_MEM_latch_out, dest4_RrAg_MEM_latch_out;
    wire         res1_ld_out_RrAg_MEM_latch_out, res2_ld_out_RrAg_MEM_latch_out, res3_ld_out_RrAg_MEM_latch_out, res4_ld_out_RrAg_MEM_latch_out;
    wire [31:0]  rep_num_RrAg_MEM_latch_out;
    wire [4:0]   aluk_RrAg_MEM_latch_out;
    wire [2:0]   mux_adder_RrAg_MEM_latch_out;
    wire         mux_and_int_RrAg_MEM_latch_out, mux_shift_RrAg_MEM_latch_out;
    wire [36:0]  p_op_RrAg_MEM_latch_out;
    wire [17:0]  fmask_RrAg_MEM_latch_out;
    wire [15:0]  CS_out_RrAg_MEM_latch_out;
    wire [1:0]   conditionals_RrAg_MEM_latch_out;
    wire         is_br_RrAg_MEM_latch_out, is_fp_RrAg_MEM_latch_out;
    wire [47:0]  imm_RrAg_MEM_latch_out;
    wire [1:0]   mem1_rw_RrAg_MEM_latch_out, mem2_rw_RrAg_MEM_latch_out;
    wire [31:0]  eip_RrAg_MEM_latch_out;
    wire         IE_RrAg_MEM_latch_out;
    wire [3:0]   IE_type_RrAg_MEM_latch_out;
    wire [31:0]  BR_pred_target_RrAg_MEM_latch_out;
    wire         BR_pred_T_NT_RrAg_MEM_latch_out;
    
    rrag r1 ( //TODO
        //inputs
        .valid_in(), .reg_addr1(), .reg_addr2(), .reg_addr3(), .reg_addr4(), .seg_addr1(), .seg_addr2(), .seg_addr3(), .seg_addr4(),
        .opsize_in(), .addressingmode(), .op1_in(), .op2_in(), .op3_in(), .op4_in(),
        .res1_ld_in(), .res2_ld_in(), .res3_ld_in(), .res4_ld_in(),
        .dest1_in(), .dest2_in(), .dest3_in(), .dest4_in(),
        .disp(), .reg3_shfamnt(), .usereg2(), .usereg3(), .rep(),
        .clr(), .clk(),
        .lim_init5(), .lim_init4(), .lim_init3(), .lim_init2(), .lim_init1(), .lim_init0(),
        .aluk_in(), .mux_adder_in(), .mux_and_int_in(), .mux_shift_in(),
        .p_op_in(), .fmask_in(), .conditionals_in(), .is_br_in(), .is_fp_in(),
        .imm_in(), .mem1_rw_in(), .mem2_rw_in(), .eip_in(), .IE_in(), .IE_type_in(),
        .BR_pred_target_in(), .BR_pred_T_NT_in(),
        .wb_data1(), .wb_data2(), .wb_data3(), .wb_data4(),
        .wb_segdata1(), .wb_segdata2(), .wb_segdata3(), .wb_segdata4(),
        .wb_addr1(), .wb_addr2(), .wb_addr3(), .wb_addr4(),
        .wb_segaddr1(), .wb_segaddr2(), .wb_segaddr3(), .wb_segaddr4(),
        .wb_opsize(), .wb_regld(), .wb_segld(), .wb_inst_ptcid(),
        .fwd_stall(),

        //outputs
        .valid_out(valid_RrAg_MEM_latch_in), .stall(stall_RrAg_MEM_latch_in), .opsize_out(opsize_RrAg_MEM_latch_in),
        .mem_addr1(mem_addr1_RrAg_MEM_latch_in), .mem_addr2(mem_addr2_RrAg_MEM_latch_in), .mem_addr1_end(mem_addr1_end_RrAg_MEM_latch_in), .mem_addr2_end(mem_addr2_end_RrAg_MEM_latch_in),
        .reg1(reg1_RrAg_MEM_latch_in), .reg2(reg2_RrAg_MEM_latch_in), .reg3(reg3_RrAg_MEM_latch_in), .reg4(reg4_RrAg_MEM_latch_in),
        .ptc_r1(ptc_r1_RrAg_MEM_latch_in), .ptc_r2(ptc_r2_RrAg_MEM_latch_in), .ptc_r3(ptc_r3_RrAg_MEM_latch_in), .ptc_r4(ptc_r4_RrAg_MEM_latch_in),
        .reg1_orig(reg1_orig_RrAg_MEM_latch_in), .reg2_orig(reg2_orig_RrAg_MEM_latch_in), .reg3_orig(reg3_orig_RrAg_MEM_latch_in), .reg4_orig(reg4_orig_RrAg_MEM_latch_in),
        .seg1(seg1_RrAg_MEM_latch_in), .seg2(seg2_RrAg_MEM_latch_in), .seg3(seg3_RrAg_MEM_latch_in), .seg4(seg4_RrAg_MEM_latch_in),
        .ptc_s1(ptc_s1_RrAg_MEM_latch_in), .ptc_s2(ptc_s2_RrAg_MEM_latch_in), .ptc_s3(ptc_s3_RrAg_MEM_latch_in), .ptc_s4(ptc_s4_RrAg_MEM_latch_in),
        .seg1_orig(seg1_orig_RrAg_MEM_latch_in), .seg2_orig(seg2_orig_RrAg_MEM_latch_in), .seg3_orig(seg3_orig_RrAg_MEM_latch_in), .seg4_orig(seg4_orig_RrAg_MEM_latch_in),
        .inst_ptcid(inst_ptcid_RrAg_MEM_latch_in),
        .op1_out(op1_out_RrAg_MEM_latch_in), .op2_out(op2_out_RrAg_MEM_latch_in), .op3_out(op3_out_RrAg_MEM_latch_in), .op4_out(op4_out_RrAg_MEM_latch_in),
        .dest1_out(dest1_out_RrAg_MEM_latch_in), .dest2_out(dest2_out_RrAg_MEM_latch_in), .dest3_out(dest3_out_RrAg_MEM_latch_in), .dest4_out(dest4_out_RrAg_MEM_latch_in),
        .res1_ld_out(res1_ld_out_RrAg_MEM_latch_in), .res2_ld_out(res2_ld_out_RrAg_MEM_latch_in), 
        .res3_ld_out(res3_ld_out_RrAg_MEM_latch_in), .res4_ld_out(res4_ld_out_RrAg_MEM_latch_in),
        .rep_num(rep_num_RrAg_MEM_latch_in),
        .aluk_out(aluk_out_RrAg_MEM_latch_in),
        .mux_adder_out(mux_adder_out_RrAg_MEM_latch_in),
        .mux_and_int_out(mux_and_int_out_RrAg_MEM_latch_in), .mux_shift_out(mux_shift_out_RrAg_MEM_latch_in),
        .p_op_out(p_op_out_RrAg_MEM_latch_in),
        .fmask_out(fmask_out_RrAg_MEM_latch_in),
        .conditionals_out(conditionals_out_RrAg_MEM_latch_in),
        .is_br_out(is_br_out_RrAg_MEM_latch_in), .is_fp_out(is_fp_out_RrAg_MEM_latch_in),
        .imm_out(imm_out_RrAg_MEM_latch_in),
        .mem1_rw_out(mem1_rw_out_RrAg_MEM_latch_in), .mem2_rw_out(mem2_rw_out_RrAg_MEM_latch_in),
        .eip_out(eip_out_RrAg_MEM_latch_in),
        .IE_out(IE_out_RrAg_MEM_latch_in),
        .IE_type_out(IE_type_out_RrAg_MEM_latch_in),
        .BR_pred_target_out(BR_pred_target_out_RrAg_MEM_latch_in),
        .BR_pred_T_NT_out(BR_pred_T_NT_out_RrAg_MEM_latch_in)
    );

    RrAg_MEM_latch q4(
        //inputs
        .valid_in(valid_RrAg_MEM_latch_in), .stall(stall_RrAg_MEM_latch_in), .opsize_in(opsize_RrAg_MEM_latch_in),
        .mem_addr1(mem_addr1_RrAg_MEM_latch_in), .mem_addr2(mem_addr2_RrAg_MEM_latch_in), .mem_addr1_end(mem_addr1_end_RrAg_MEM_latch_in), .mem_addr2_end(mem_addr2_end_RrAg_MEM_latch_in),
        .reg1(reg1_RrAg_MEM_latch_in), .reg2(reg2_RrAg_MEM_latch_in), .reg3(reg3_RrAg_MEM_latch_in), .reg4(reg4_RrAg_MEM_latch_in),
        .ptc_r1(ptc_r1_RrAg_MEM_latch_in), .ptc_r2(ptc_r2_RrAg_MEM_latch_in), .ptc_r3(ptc_r3_RrAg_MEM_latch_in), .ptc_r4(ptc_r4_RrAg_MEM_latch_in),
        .reg1_orig(reg1_orig_RrAg_MEM_latch_in), .reg2_orig(reg2_orig_RrAg_MEM_latch_in), .reg3_orig(reg3_orig_RrAg_MEM_latch_in), .reg4_orig(reg4_orig_RrAg_MEM_latch_in),
        .seg1(seg1_RrAg_MEM_latch_in), .seg2(seg2_RrAg_MEM_latch_in), .seg3(seg3_RrAg_MEM_latch_in), .seg4(seg4_RrAg_MEM_latch_in),
        .ptc_s1(ptc_s1_RrAg_MEM_latch_in), .ptc_s2(ptc_s2_RrAg_MEM_latch_in), .ptc_s3(ptc_s3_RrAg_MEM_latch_in), .ptc_s4(ptc_s4_RrAg_MEM_latch_in),
        .seg1_orig(seg1_orig_RrAg_MEM_latch_in), .seg2_orig(seg2_orig_RrAg_MEM_latch_in), .seg3_orig(seg3_orig_RrAg_MEM_latch_in), .seg4_orig(seg4_orig_RrAg_MEM_latch_in),
        .inst_ptcid(inst_ptcid_RrAg_MEM_latch_in),
        .op1_sel(op1_out_RrAg_MEM_latch_in), .op2_sel(op2_out_RrAg_MEM_latch_in), .op3_sel(op3_out_RrAg_MEM_latch_in), .op4_sel(op4_out_RrAg_MEM_latch_in),
        .dest1_sel(dest1_out_RrAg_MEM_latch_in), .dest2_sel(dest2_out_RrAg_MEM_latch_in), .dest3_sel(dest3_out_RrAg_MEM_latch_in), .dest4_sel(dest4_out_RrAg_MEM_latch_in),
        .res1_ld_in(res1_ld_out_RrAg_MEM_latch_in), .res2_ld_in(res2_ld_out_RrAg_MEM_latch_in),
        .res3_ld_in(res3_ld_out_RrAg_MEM_latch_in), .res4_ld_in(res4_ld_out_RrAg_MEM_latch_in),
        .rep_num(rep_num_RrAg_MEM_latch_in),
        .aluk_in(aluk_out_RrAg_MEM_latch_in), .mux_adder_in(mux_adder_out_RrAg_MEM_latch_in),
        .mux_and_int_in(mux_and_int_out_RrAg_MEM_latch_in), .mux_shift_in(mux_shift_out_RrAg_MEM_latch_in),
        .p_op_in(p_op_out_RrAg_MEM_latch_in), .fmask_in(fmask_out_RrAg_MEM_latch_in),
        .conditionals_in(conditionals_out_RrAg_MEM_latch_in), .is_br_in(is_br_out_RrAg_MEM_latch_in),
        .is_fp_in(is_fp_out_RrAg_MEM_latch_in),
        .imm(imm_out_RrAg_MEM_latch_in), .mem1_rw(mem1_rw_out_RrAg_MEM_latch_in), .mem2_rw(mem2_rw_out_RrAg_MEM_latch_in),
        .eip_in(eip_out_RrAg_MEM_latch_in), .IE_in(IE_out_RrAg_MEM_latch_in), .IE_type_in(IE_type_out_RrAg_MEM_latch_in),
        .BR_pred_target_in(BR_pred_target_out_RrAg_MEM_latch_in), .BR_pred_T_NT_in(BR_pred_T_NT_out_RrAg_MEM_latch_in),
        .clk(clk),
        //outputs

        .valid_out(valid_RrAg_MEM_latch_out), .stall(stall_RrAg_MEM_latch_out), .opsize_out(opsize_RrAg_MEM_latch_out),
        .mem_addr1(mem_addr1_RrAg_MEM_latch_out), .mem_addr2(mem_addr2_RrAg_MEM_latch_out), .mem_addr1_end(mem_addr1_end_RrAg_MEM_latch_out), .mem_addr2_end(mem_addr2_end_RrAg_MEM_latch_out),
        .reg1(reg1_RrAg_MEM_latch_out), .reg2(reg2_RrAg_MEM_latch_out), .reg3(reg3_RrAg_MEM_latch_out), .reg4(reg4_RrAg_MEM_latch_out),
        .ptc_r1(ptc_r1_RrAg_MEM_latch_out), .ptc_r2(ptc_r2_RrAg_MEM_latch_out), .ptc_r3(ptc_r3_RrAg_MEM_latch_out), .ptc_r4(ptc_r4_RrAg_MEM_latch_out),
        .reg1_orig(reg1_orig_RrAg_MEM_latch_out), .reg2_orig(reg2_orig_RrAg_MEM_latch_out), .reg3_orig(reg3_orig_RrAg_MEM_latch_out), .reg4_orig(reg4_orig_RrAg_MEM_latch_out),
        .seg1(seg1_RrAg_MEM_latch_out), .seg2(seg2_RrAg_MEM_latch_out), .seg3(seg3_RrAg_MEM_latch_out), .seg4(seg4_RrAg_MEM_latch_out),
        .ptc_s1(ptc_s1_RrAg_MEM_latch_out), .ptc_s2(ptc_s2_RrAg_MEM_latch_out), .ptc_s3(ptc_s3_RrAg_MEM_latch_out), .ptc_s4(ptc_s4_RrAg_MEM_latch_out),
        .seg1_orig(seg1_orig_RrAg_MEM_latch_out), .seg2_orig(seg2_orig_RrAg_MEM_latch_out), .seg3_orig(seg3_orig_RrAg_MEM_latch_out), .seg4_orig(seg4_orig_RrAg_MEM_latch_out),
        .inst_ptcid(inst_ptcid_RrAg_MEM_latch_out),
        .op1_sel(op1_RrAg_MEM_latch_out), .op2_sel(op2_RrAg_MEM_latch_out), .op3_sel(op3_RrAg_MEM_latch_out), .op4_sel(op4_RrAg_MEM_latch_out),
        .dest1_sel(dest1_RrAg_MEM_latch_out), .dest2_sel(dest2_RrAg_MEM_latch_out), .dest3_sel(dest3_RrAg_MEM_latch_out), .dest4_sel(dest4_RrAg_MEM_latch_out),
        .res1_ld_in(res1_ld_out_RrAg_MEM_latch_out), .res2_ld_in(res2_ld_out_RrAg_MEM_latch_out),
        .res3_ld_in(res3_ld_out_RrAg_MEM_latch_out), .res4_ld_in(res4_ld_out_RrAg_MEM_latch_out),
        .rep_num(rep_num_RrAg_MEM_latch_out),
        .aluk_in(aluk_RrAg_MEM_latch_out), .mux_adder_in(mux_adder_RrAg_MEM_latch_out),
        .mux_and_int_in(mux_and_int_RrAg_MEM_latch_out), .mux_shift_in(mux_shift_RrAg_MEM_latch_out),
        .p_op_in(p_op_RrAg_MEM_latch_out), .fmask_in(fmask_RrAg_MEM_latch_out),
        .conditionals_in(conditionals_RrAg_MEM_latch_out), .is_br_in(is_br_RrAg_MEM_latch_out),
        .is_fp_in(is_fp_RrAg_MEM_latch_out),
        .imm(imm_RrAg_MEM_latch_out), .mem1_rw(mem1_rw_RrAg_MEM_latch_out), .mem2_rw(mem2_rw_RrAg_MEM_latch_out),
        .eip_in(eip_RrAg_MEM_latch_out), .IE_in(IE_RrAg_MEM_latch_out), .IE_type_in(IE_type_RrAg_MEM_latch_out),
        .BR_pred_target_in(BR_pred_target_RrAg_MEM_latch_out), .BR_pred_T_NT_in(BR_pred_T_NT_RrAg_MEM_latch_out)
    );


    mem m1 (
        .valid_in(valid_RrAg_MEM_latch_out),
        .opsize_in(opsize_RrAg_MEM_latch_out),
        .mem_addr1(mem_addr1_RrAg_MEM_latch_out),
        .mem_addr2(mem_addr2_RrAg_MEM_latch_out),
        .mem_addr1_end(mem_addr1_end_RrAg_MEM_latch_out),
        .mem_addr2_end(mem_addr2_end_RrAg_MEM_latch_out),
        .reg1(reg1_RrAg_MEM_latch_out),
        .reg2(reg2_RrAg_MEM_latch_out),
        .reg3(reg3_RrAg_MEM_latch_out),
        .reg4(reg4_RrAg_MEM_latch_out),
        .ptc_r1(ptc_r1_RrAg_MEM_latch_out),
        .ptc_r2(ptc_r2_RrAg_MEM_latch_out),
        .ptc_r3(ptc_r3_RrAg_MEM_latch_out),
        .ptc_r4(ptc_r4_RrAg_MEM_latch_out),
        .reg1_orig(reg1_orig_RrAg_MEM_latch_out),
        .reg2_orig(reg2_orig_RrAg_MEM_latch_out),
        .reg3_orig(reg3_orig_RrAg_MEM_latch_out),
        .reg4_orig(reg4_orig_RrAg_MEM_latch_out),
        .seg1(seg1_RrAg_MEM_latch_out),
        .seg2(seg2_RrAg_MEM_latch_out),
        .seg3(seg3_RrAg_MEM_latch_out),
        .seg4(seg4_RrAg_MEM_latch_out),
        .ptc_s1(ptc_s1_RrAg_MEM_latch_out),
        .ptc_s2(ptc_s2_RrAg_MEM_latch_out),
        .ptc_s3(ptc_s3_RrAg_MEM_latch_out),
        .ptc_s4(ptc_s4_RrAg_MEM_latch_out),
        .seg1_orig(seg1_orig_RrAg_MEM_latch_out),
        .seg2_orig(seg2_orig_RrAg_MEM_latch_out),
        .seg3_orig(seg3_orig_RrAg_MEM_latch_out),
        .seg4_orig(seg4_orig_RrAg_MEM_latch_out),
        .inst_ptcid(inst_ptcid_RrAg_MEM_latch_out),
        .op1_sel(op1_RrAg_MEM_latch_out),
        .op2_sel(op2_RrAg_MEM_latch_out),
        .op3_sel(op3_RrAg_MEM_latch_out),
        .op4_sel(op4_RrAg_MEM_latch_out),
        .dest1_sel(dest1_RrAg_MEM_latch_out),
        .dest2_sel(dest2_RrAg_MEM_latch_out),
        .dest3_sel(dest3_RrAg_MEM_latch_out),
        .dest4_sel(dest4_RrAg_MEM_latch_out),
        .res1_ld_in(res1_ld_out_RrAg_MEM_latch_out), .res2_ld_in(res2_ld_out_RrAg_MEM_latch_out),
        .res3_ld_in(res3_ld_out_RrAg_MEM_latch_out), .res4_ld_in(res4_ld_out_RrAg_MEM_latch_out),
        .rep_num(rep_num_RrAg_MEM_latch_out),
        .VP_in(VP), .PF_in(PF),
        .entry_v_in(entry_v), .entry_P_in(entry_P), .entry_RW_in(entry_RW), .entry_PCD_in(entry_PCD),
        .aluk_in(aluk_RrAg_MEM_latch_out), .mux_adder_in(mux_adder_RrAg_MEM_latch_out), 
        .mux_and_int_in(mux_and_int_RrAg_MEM_latch_out), .mux_shift_in(mux_shift_RrAg_MEM_latch_out),
        .p_op_in(p_op_RrAg_MEM_latch_out), .fmask_in(fmask_RrAg_MEM_latch_out),
        .CS_in(CS_out_RrAg_MEM_latch_out),
        .conditionals_in(conditionals_RrAg_MEM_latch_out), .is_br_in(is_br_RrAg_MEM_latch_out), 
        .is_fp_in(is_fp_RrAg_MEM_latch_out),
        .imm(imm_RrAg_MEM_latch_out), .mem1_rw(mem1_rw_RrAg_MEM_latch_out), .mem2_rw(mem2_rw_RrAg_MEM_latch_out),
        .eip_in(eip_RrAg_MEM_latch_out), .IE_in(IE_RrAg_MEM_latch_out), .IE_type_in(IE_type_RrAg_MEM_latch_out),
        .BR_pred_target_in(BR_pred_target_RrAg_MEM_latch_out), .BR_pred_T_NT_in(BR_pred_T_NT_RrAg_MEM_latch_out),
        .clr(/*TODO*/), .clk(clk),
        //outputs
        .valid_out(valid_MEM_EX_latch_in),
        .eip_out(EIP_MEM_EX_latch_in),
        .IE_out(IE_MEM_EX_latch_in),
        .IE_type_out(IE_type_MEM_EX_latch_in),
        .BR_pred_target_out(BR_pred_target_MEM_EX_latch_in),
        .BR_pred_T_NT_out(BR_pred_T_NT_MEM_EX_latch_in),
        .opsize_out(opsize_MEM_EX_latch_in)
        .set_out(set_MEM_EX_latch_in),
        .rst_out(rst_MEM_EX_latch_in),
        .res1_ld_out(res1_ld_MEM_EX_latch_in),
        .res2_ld_out(res2_ld_MEM_EX_latch_in),
        .res3_ld_out(res3_ld_MEM_EX_latch_in),
        .res4_ld_out(res4_ld_MEM_EX_latch_in),
        .op1_val(op1_MEM_EX_latch_in),
        .op2_val(op2_MEM_EX_latch_in),
        .op3_val(op3_MEM_EX_latch_in),
        .op4_val(op4_MEM_EX_latch_in),
        .op1_ptcinfo(op1_ptcinfo_MEM_EX_latch_in),
        .op2_ptcinfo(op2_ptcinfo_MEM_EX_latch_in),
        .op3_ptcinfo(op3_ptcinfo_MEM_EX_latch_in),
        .op4_ptcinfo(op4_ptcinfo_MEM_EX_latch_in),
        .dest1_addr(dest1_addr_MEM_EX_latch_in),
        .dest2_addr(dest2_addr_MEM_EX_latch_in),
        .dest3_addr(dest3_addr_MEM_EX_latch_in),
        .dest4_addr(dest4_addr_MEM_EX_latch_in),
        .dest1_is_reg(res1_is_reg_MEM_EX_latch_in),
        .dest2_is_reg(res2_is_reg_MEM_EX_latch_in),
        .dest3_is_reg(res3_is_reg_MEM_EX_latch_in),
        .dest4_is_reg(res4_is_reg_MEM_EX_latch_in),
        .dest1_is_seg(res1_is_seg_MEM_EX_latch_in),
        .dest2_is_seg(res2_is_seg_MEM_EX_latch_in),
        .dest3_is_seg(res3_is_seg_MEM_EX_latch_in),
        .dest4_is_seg(res4_is_seg_MEM_EX_latch_in),
        .dest1_is_mem(res1_is_mem_MEM_EX_latch_in), .dest2_is_mem(res2_is_mem_MEM_EX_latch_in), 
        .dest3_is_mem(res3_is_mem_MEM_EX_latch_in), .dest4_is_mem(res4_is_mem_MEM_EX_latch_in),
        .aluk_out(aluk_MEM_EX_latch_in), .mux_adder_out(MUX_ADDER_IMM_MEM_EX_latch_in), 
        .mux_and_int_out(MUX_AND_INT_MEM_EX_latch_in), .mux_shift_out(MUX_SHIFT_MEM_EX_latch_in),
        .p_op_out(P_OP_MEM_EX_latch_in), .fmask_out(FMASK_MEM_EX_latch_in), .conditionals_out(conditionals_MEM_EX_latch_in), .is_br_out(isBR_MEM_EX_latch_in), .is_fp_out(is_fp_MEM_EX_latch_in),
        .CS_out(CS_MEM_EX_latch_in)
    );        
        
    ///////////////////////////////////////////////////////////
    //     Outputs from EX that go into EX_WB_latch:        //  
    //////////////////////////////////////////////////////////

    wire valid_MEM_EX_latch_in;
    wire [31:0] EIP_MEM_EX_latch_in;
    wire IE_MEM_EX_latch_in;
    wire [3:0] IE_type_MEM_EX_latch_in;
    wire [31:0] BR_pred_target_MEM_EX_latch_in;
    wire BR_pred_T_NT_MEM_EX_latch_in;

    wire res1_ld_MEM_EX_latch_in, res2_ld_MEM_EX_latch_in, res3_ld_MEM_EX_latch_in, res4_ld_MEM_EX_latch_in;
    wire [63:0] op1_MEM_EX_latch_in, op2_MEM_EX_latch_in, op3_MEM_EX_latch_in, op4_MEM_EX_latch_in;
    wire [127:0] op1_ptcinfo_MEM_EX_latch_in, op2_ptcinfo_MEM_EX_latch_in, op3_ptcinfo_MEM_EX_latch_in, op4_ptcinfo_MEM_EX_latch_in;
    wire [31:0] dest1_addr_MEM_EX_latch_in, dest2_addr_MEM_EX_latch_in, dest3_addr_MEM_EX_latch_in, dest4_addr_MEM_EX_latch_in;
    wire res1_is_reg_MEM_EX_latch_in, res2_is_reg_MEM_EX_latch_in, res3_is_reg_MEM_EX_latch_in, res4_is_reg_MEM_EX_latch_in;
    wire res1_is_seg_MEM_EX_latch_in, res2_is_seg_MEM_EX_latch_in, res3_is_seg_MEM_EX_latch_in, res4_is_seg_MEM_EX_latch_in;
    wire res1_is_mem_MEM_EX_latch_in, res2_is_mem_MEM_EX_latch_in, res3_is_mem_MEM_EX_latch_in, res4_is_mem_MEM_EX_latch_in;
    wire [1:0] opsize_MEM_EX_latch_in;

    wire [4:0] aluk_MEM_EX_latch_in;
    wire [2:0] MUX_ADDER_IMM_MEM_EX_latch_in;
    wire MUX_AND_INT_MEM_EX_latch_in, MUX_SHIFT_MEM_EX_latch_in;

    wire [34:0] P_OP_MEM_EX_latch_in;
    wire [16:0] FMASK_MEM_EX_latch_in;
    wire [1:0] conditionals_MEM_EX_latch_in;

    wire isBR_MEM_EX_latch_in, is_fp_MEM_EX_latch_in;
    wire [15:0] CS_MEM_EX_latch_in;

    ///////////////////////////////////////////////////////////
    //     Outputs from EX_WB_latch that go into WB:        //  
    //////////////////////////////////////////////////////////

    wire valid_MEM_EX_latch_out;
    wire [31:0] EIP_MEM_EX_latch_out;
    wire IE_MEM_EX_latch_out;
    wire [3:0] IE_type_MEM_EX_latch_out;
    wire [31:0] BR_pred_target_MEM_EX_latch_out;
    wire BR_pred_T_NT_MEM_EX_latch_out;

    wire res1_ld_MEM_EX_latch_out, res2_ld_MEM_EX_latch_out, res3_ld_MEM_EX_latch_out, res4_ld_MEM_EX_latch_out;
    wire [63:0] op1_MEM_EX_latch_out, op2_MEM_EX_latch_out, op3_MEM_EX_latch_out, op4_MEM_EX_latch_out;
    wire [127:0] op1_ptcinfo_MEM_EX_latch_out, op2_ptcinfo_MEM_EX_latch_out, op3_ptcinfo_MEM_EX_latch_out, op4_ptcinfo_MEM_EX_latch_out;
    wire [31:0] dest1_addr_MEM_EX_latch_out, dest2_addr_MEM_EX_latch_out, dest3_addr_MEM_EX_latch_out, dest4_addr_MEM_EX_latch_out;
    wire res1_is_reg_MEM_EX_latch_out, res2_is_reg_MEM_EX_latch_out, res3_is_reg_MEM_EX_latch_out, res4_is_reg_MEM_EX_latch_out;
    wire res1_is_seg_MEM_EX_latch_out, res2_is_seg_MEM_EX_latch_out, res3_is_seg_MEM_EX_latch_out, res4_is_seg_MEM_EX_latch_out;
    wire res1_is_mem_MEM_EX_latch_out, res2_is_mem_MEM_EX_latch_out, res3_is_mem_MEM_EX_latch_out, res4_is_mem_MEM_EX_latch_out;
    wire [1:0] opsize_MEM_EX_latch_out;

    wire [4:0] aluk_MEM_EX_latch_out;
    wire [2:0] MUX_ADDER_IMM_MEM_EX_latch_out;
    wire MUX_AND_INT_MEM_EX_latch_out, MUX_SHIFT_MEM_EX_latch_out;
    wire [34:0] P_OP_MEM_EX_latch_out;
    wire [16:0] FMASK_MEM_EX_latch_out;
    wire [1:0] conditionals_MEM_EX_latch_out;

    wire isBR_MEM_EX_latch_out, is_fp_MEM_EX_latch_out;
    wire [15:0] CS_MEM_EX_latch_out;

    //queued latches between MEM and EX - 8

    integer m_size, n_size;

    wire [m_size-1:0] m_din;
    wire [n_size-1:0] n_din;

    MEM_EX_Queued_Latches #(.M_WIDTH(/*TODO*/), .N_WIDTH(/*TODO*/), .Q_LENGTH(8)) q5 (
        .m_din(/*TODO*/), .n_din(/*TODO*/), .new_m_vector(/*TODO*/), .wr(/*TODO*/), .rd(/*TODO*/), 
        .modify_vector(/*TODO*/), .clr(/*TODO*/), .clk(clk), .full(/*TODO*/), .empty(/*TODO*/), .old_m_vector(/*TODO*/), .dout(/*TODO*/)
    );

    execute_TOP e1 (
        .clk(clk),
        .valid_in(valid_MEM_EX_latch_out),
        .EIP_in(EIP_MEM_EX_latch_out),
        .IE_in(IE_MEM_EX_latch_out),  
        .IE_type_in(IE_type_MEM_EX_latch_out),
        .BR_pred_target_in(BR_pred_target_MEM_EX_latch_out),     
        .BR_pred_T_NT_in(BR_pred_T_NT_MEM_EX_latch_out),        
        .set(), .rst(), //TODO

        .res1_ld_in(res1_ld_MEM_EX_latch_out), .res2_ld_in(res2_ld_MEM_EX_latch_out),
        .res3_ld_in(res3_ld_MEM_EX_latch_out), .res4_ld_in(res4_ld_MEM_EX_latch_out),
        .op1(op1_MEM_EX_latch_out), .op2(op2_MEM_EX_latch_out),
        .op3(op2_MEM_EX_latch_out), .op4(op4_MEM_EX_latch_out),
        .op1_ptcinfo(op1_ptcinfo_MEM_EX_latch_out), .op2_ptcinfo(op2_ptcinfo_MEM_EX_latch_out),
        .op3_ptcinfo(op3_ptcinfo_MEM_EX_latch_out), .op4_ptcinfo(op4_ptcinfo_MEM_EX_latch_out),
        .dest1_addr(dest1_addr_MEM_EX_latch_out), .dest2_addr(dest2_addr_MEM_EX_latch_out), 
        .dest3_addr(dest3_addr_MEM_EX_latch_out), .dest4_addr(dest4_addr_MEM_EX_latch_out),
        .res1_is_reg_in(res1_is_reg_MEM_EX_latch_out), .res2_is_reg_in(res2_is_reg_MEM_EX_latch_out),
        .res3_is_reg_in(res3_is_reg_MEM_EX_latch_out), .res4_is_reg_in(res4_is_reg_MEM_EX_latch_out),
        .res1_is_seg_in(res1_is_seg_MEM_EX_latch_out), .res2_is_seg_in(res2_is_seg_MEM_EX_latch_out),
        .res3_is_seg_in(res3_is_seg_MEM_EX_latch_out), .res4_is_seg_in(res4_is_seg_MEM_EX_latch_out),
        .res1_is_mem_in(res1_is_mem_MEM_EX_latch_out), .res2_is_mem_in(res2_is_mem_MEM_EX_latch_out), 
        .res3_is_mem_in(res3_is_mem_MEM_EX_latch_out), .res4_is_mem_in(res4_is_mem_MEM_EX_latch_out),
        .opsize_in(opsize_MEM_EX_latch_out),
        
        .aluk(aluk_MEM_EX_latch_out),
        .MUX_ADDER_IMM(MUX_ADDER_IMM_MEM_EX_latch_out),
        .MUX_AND_INT(MUX_AND_INT_MEM_EX_latch_out),
        .MUX_SHIFT(MUX_SHIFT_MEM_EX_latch_out),
        .P_OP(P_OP_MEM_EX_latch_out),
        .FMASK(FMASK_MEM_EX_latch_out),
        .conditionals(conditionals_MEM_EX_latch_out),    
        .isBR(isBR_MEM_EX_latch_out),
        .is_fp(is_fp_MEM_EX_latch_out), 
        .CS(CS_MEM_EX_latch_out),
        
        //outputs:
        .valid_out(),
        .EIP_out(),
        .IE_out(),
        .IE_type_out(),
        .BR_pred_target_out(),
        .BR_pred_T_NT_out(),
        
        .eflags(),
        .CS_out(), 
        
        .res1_wb(), .res2_wb(), .res3_wb(), .res4_wb(),
        .res1(), .res2(), res3(), .res4(),
        .res1_is_reg_out(), .res2_is_reg_out(), .res3_is_reg_out(), .res4_is_reg_out(), 
        .res1_is_seg_out(), .res2_is_seg_out(), .res3_is_seg_out(), .res4_is_seg_out(), 
        .res1_is_mem_out(), .res2_is_mem_out(), .res3_is_mem_out(), .res4_is_mem_out(),
        .res1_dest(), .res2_dest(), .res3_dest(), .res4_dest(), 
        .ressize(), 

        .BR_valid(), 
        .BR_taken(),
        .BR_correct(), 
        .BR_FIP(), 
        .BR_FIP_p1()
    );


endmodule

