module bp_gshare (
    input [31:0] eip

);


endmodule