module DMA(
    input clk,
    input set, rst,
    
    //DES
    output reg read_d,
    
    input full_d,
    input [14:0] pAdr_d,
    input [16*8-1:0] data_d,
    input [3:0]return_d,
    input [3:0] dest_d,
    input rw_d,
    input [15:0] size_d,

    //S
    output reg valid_s,
    output reg [14:0] pAdr_s,
    output reg [16*8-1:0] data_s,
    output reg [3:0] dest_s,
    output reg [3:0]return_s,
    output reg rw_s,
    output reg [15:0] size_s,

    input full_block_s,
    input free_block_s,

    //DISC
    input [127:0] data_disc,
    input finished_disc,
    output reg [32:0] adr_disc,
    output reg read_disc,

    //KEYBOARD
    input [7:0] data_kb,
    output reg read_kb,

    //CORE
    output wire interrupt_core
);
//ADDRESS_LIST
//readCHAR: x1000
//Disc Source: x1010
//Memory destination: x1020
//Disc size: x1030
//Initialize: x1040
//ClearInterrupt x1050
reg interrupt;
assign interrupt_core = interrupt;

reg[31:0] discSource;
reg[14:0] memDest;
reg[11:0] discSize;
reg inUse;
wire[127:0] ldSER;

reg [127:0] discBuffer;
reg[3:0] state;

concat_io a(discSize[3:0], data_d, discBuffer[127:0], ldSER);
reg[4095:0] upCnt;
always @(posedge clk) begin
    if(!rst) begin
        inUse = 0;
        memDest = 0;
        discSource = 0;
        discSize = 0;
        valid_s = 0;
        read_d = 0;
        interrupt = 0;
        discBuffer = 0;
        upCnt = 0;
        state = 0;
        adr_disc = 33'h1_0000_0000;

    end
    else begin 
        case(state)
            4'b0000: begin
                read_kb = 0;
                read_d = 0;
                valid_s = 0;
                if(full_d) begin 
                    case (pAdr_d[6:4])
                        3'b000: begin                          
                                read_kb = 1;
                                state = 1;
                        end

                        3'b001: begin
                            discSource = data_d[31:0];
                            read_d = 1;
                        end

                        3'b010: begin
                            memDest = data_d[14:0];
                            read_d = 1;
                        end

                        3'b011: begin
                            discSize = data_d[11:0];
                            read_d = 1;
                        end

                        3'b100: begin
                                state = 4;
                                read_d = 1;
                                adr_disc = {1'b0,discSource};
                                upCnt = 0;
                            
                        end

                        3'b101: begin
                            interrupt = 0;
                            read_d = 1'b1;
                        end
                        default: begin
                            read_d = 1'b1;
                        end
                    endcase
                end
            else begin
                read_kb = 0;
                read_d = 0;
                valid_s = 0;
            end
            end
            
            4'b0001:begin
                read_kb = 0;
                read_d = 0;
                valid_s = 0;
                if(free_block_s) begin
                    valid_s=1;
                    pAdr_s = pAdr_d;
                    data_s = {120'd0, data_kb};
                    return_s = 4'b1100;
                    dest_s = return_d;
                    rw_s = 1'b1;
                    size_s = 16'h8000;
                    state = 0;
                end
            end

            4'b0011: begin
                valid_s = 0;
                read_d = 0;
                read_disc = 0;
                if(free_block_s) begin
                    valid_s=1;
                    pAdr_s = pAdr_d;
                    data_s = {120'd0, data_kb};
                    return_s = 4'b1100;
                    dest_s = return_d;
                    rw_s =  1'b1;
                    size_s = 16'h8000;
                    state = 4'b0100;
                end
            end

            4'b0100: begin
                valid_s = 0;
                read_d = 0;
                read_disc = 0;
                inUse = 1;
                read_d = 1;
                adr_disc = {1'b0,discSource};
                upCnt = 0;
                if(finished_disc)begin
                    discBuffer = data_disc;
                    read_disc = 1;
                    if(discSize > 16) state = 4'b0110;
                  else state = 4'b0111;
                end
            end

            4'b0110: begin
                valid_s = 0;
                read_d = 0;
                read_disc = 0;
                if(free_block_s) begin 
                    if(pAdr_d[6:4] == 3'b000)begin
                        valid_s=1;
                        pAdr_s = pAdr_d;
                        data_s = {120'd0, data_kb};
                        return_s = 4'b1100;
                        dest_s = return_d;
                        rw_s =  1'b1;
                        size_s = 16'h8000;
                        read_d = 1;
                    end
                    else begin
                        valid_s <=1 ;
                        pAdr_s <= memDest;
                        data_s <= discBuffer;
                        return_s <= 4'b1100;
                        dest_s <= {2'b10, memDest[1:0]};
                        rw_s <= 1'b1;
                        size_s <= 16'h8000;
                        upCnt <= upCnt + 127;
                        discSource <= discSource + 32'h0010;
                        memDest <= memDest + 16;
                        if(discSize > 16) state <= 4'b0100;
                        else state <= 4'b0111;
                        discSize <= discSize - 16;
                    end
                end
            end

        4'b0111: begin 
            valid_s = 0;
                read_d = 0;
                read_disc = 0;
            if(free_block_s) begin
                valid_s =1 ;
                pAdr_s = memDest;
                data_s = discBuffer[  127 : 0];
                return_s = 4'b1100;
                dest_s = {2'b10, memDest[1:0]};
                rw_s = 1'b0;
                size_s = 16'h1000;
                upCnt = upCnt + 127;
                discSource = discSource + 32'h0010;
                memDest = memDest + 16;
                discSize = discSize - 16;
                state = 4'b1000;
            end
        end
        4'b1000: begin
            read_kb = 0;
                read_d = 0;
                valid_s = 0;
            if(free_block_s)begin
                if(full_d) begin
                    valid_s =1 ;
                    pAdr_s = memDest;
                    data_s = ldSER;
                    return_s = 4'b1100;
                    dest_s = {2'b10, memDest[1:0]};
                    rw_s = 1'b1;
                    size_s = 16'h8000;
                    upCnt = upCnt + 127;
                    discSize = 0;
                    memDest = memDest + 16;
                    interrupt = 1;
                    state = 4'b1001;
                end
            end
        end

        4'b1001: begin
            read_kb = 0;
                read_d = 0;
                valid_s = 0;
            state = 0; 
            interrupt = 0;
            end            
        endcase
    end
end 



endmodule



module concat_io(
    input[3:0] discSize,
    input [127:0] fromMem,
    input[127:0] fromDisc, 
    output reg [127:0] toMem);

    always @(*) begin
        case(discSize)
        4'd0: toMem = fromMem;
        4'd1: toMem = {fromMem[127:8],fromDisc[7:0]};
        4'd2: toMem = {fromMem[127:16],fromDisc[15:0]};
        4'd3: toMem = {fromMem[127:24],fromDisc[23:0]};
        4'd4: toMem = {fromMem[127:32],fromDisc[31:0]};
        4'd5: toMem = {fromMem[127:40],fromDisc[39:0]};
        4'd6: toMem = {fromMem[127:48],fromDisc[47:0]};
        4'd7: toMem = {fromMem[127:56],fromDisc[55:0]};
        4'd8: toMem = {fromMem[127:64],fromDisc[63:0]};
        4'd9: toMem = {fromMem[127:72],fromDisc[71:0]};
        4'd10: toMem = {fromMem[127:80],fromDisc[79:0]};
        4'd11: toMem = {fromMem[127:88],fromDisc[87:0]};
        4'd12: toMem = {fromMem[127:96],fromDisc[95:0]};
        4'd13: toMem = {fromMem[127:104],fromDisc[103:0]};
        4'd14: toMem = {fromMem[127:112],fromDisc[111:0]};
        4'd15: toMem = {fromMem[127:120],fromDisc[119:0]};
        default: toMem = fromDisc;
        endcase
    end



endmodule
/*if(full_d) begin
            valid_s = 0;
            read_kb = 0;
            if(inUse && state == 3) begin 
                        if(free_block_s) begin
                            valid_s =1 ;
                            pAdr_s = memDest;
                            data_s = ldSER;
                            return_s = 4'b1100;
                            dest_s = {2'b10, memDest[1:0]};
                            rw_s = 1'b1;
                            size_s = 16'h8000;
                            upCnt = upCnt + 127;
                            discSize = discSize - 16;
                            memDest = memDest + 16;
                            interrupt = 1;
                        end
            end
            else begin
                $display("pAdr_d 6 - 4 0x%0h\n", pAdr_d[6:4]);
            case (pAdr_d[6:4])
                
                3'b000: begin
                    if(free_block_s) begin                        
                        read_kb = 1;
                    end 
                end

                3'b001: begin
                    discSource = inUse? discSource: data_d[31:0];
                    read_d = 1;
                end

                3'b010: begin
                    memDest = inUse? memDest:data_d[14:0];
                    read_d = 1;
                end

                3'b011: begin
                    discSize = inUse? discSize:data_d[11:0];
                    read_d = 1;
                end

                3'b100: begin
                    
                        inUse = 1;
                        state = 1;
                        read_d = 1;
                        adr_disc = {1'b0,discSource};
                        upCnt = 0;
                    
                end

                3'b101: begin
                    interrupt = 0;
                     read_d = 1'b1;
                end
                default: begin
                    read_d = 1'b1;
                end
            endcase
        end
    
        
        
        end
        else begin 
            read_kb = 0;
            read_d = 0;
            valid_s = 0;
        end

        if(free_block_s) begin
                if(pAdr_d[6:4] == 3'b000)begin
                    valid_s=1;
                    pAdr_s = pAdr_d;
                    data_s = {120'd0, data_kb};
                    return_s = 4'b1100;
                    dest_s = return_d;
                    rw_s = ~ rw_d;
                    size_s = 16'h8000;
                end
                else if(inUse) begin
                    if(state == 1 && finished_disc ) begin 
                        state = 2;
                        discBuffer = data_disc;
                    end
                    else if(state == 2) begin
                        if(discSize < 16) begin 
                            if(discSize == 0) begin
                                inUse = 0;
                                state = 0;
                                interrupt = 1;
                            end
                            else begin
                                state = 3;
                                valid_s =1 ;
                                pAdr_s = memDest;
                                data_s = discBuffer[  127 :0 ];
                                return_s = 4'b1100;
                                dest_s = {2'b10, memDest[1:0]};
                                rw_s = 1'b0;
                                size_s = 16'h8000;
                                upCnt = upCnt;
                                discSize = 0;
                                memDest = memDest;
                            end
                        end
                        else begin
                            valid_s =1 ;
                            pAdr_s = memDest;
                            data_s = discBuffer[  127 : 0];
                            return_s = 4'b1100;
                            dest_s = {2'b10, memDest[1:0]};
                            rw_s = 1'b1;
                            size_s = 16'h8000;
                            upCnt = upCnt + 127;
                            discSize = discSize - 16;
                            memDest = memDest + 16;
                            discBuffer = discBuffer >> 128;
                        end
                    end
                end
        end


    end 
    */