module skipgen_t();

endmodule